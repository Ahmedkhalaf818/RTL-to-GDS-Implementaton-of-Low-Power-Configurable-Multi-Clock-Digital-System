

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO SYS_TOP 
  PIN SI[4] 
    ANTENNAPARTIALMETALAREA 1.923 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.24963 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.498 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.39778 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.168 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.00048 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 29.46 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 141.895 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 575.66 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2781.57 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA56 ;
  END SI[4]
  PIN SI[3] 
    ANTENNAPARTIALMETALAREA 0.337 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.62097 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.432 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 2.27032 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 4.664 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 22.6262 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 31.51 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 151.756 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 649.468 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 3137.73 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 3.38649 LAYER VIA56 ;
  END SI[3]
  PIN SI[2] 
    ANTENNAPARTIALMETALAREA 2.505 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 12.0491 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.25 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3949 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 21.26 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 102.453 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 436.391 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2112.83 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 4.74109 LAYER VIA56 ;
  END SI[2]
  PIN SI[1] 
    ANTENNAPARTIALMETALAREA 1.973 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.49013 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 3.525 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.1476 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 111.382 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 542.315 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.3546 LAYER VIA34 ;
  END SI[1]
  PIN SI[0] 
    ANTENNAPARTIALMETALAREA 2.169 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 10.4329 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.017 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.5142 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 8.632 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 41.7123 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 187.01 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 909.698 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.70919 LAYER VIA45 ;
  END SI[0]
  PIN SO[4] 
    ANTENNADIFFAREA 0.537 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 8.228 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 39.7691 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 48.4448 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 233.405 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.81104 LAYER VIA34 ;
  END SO[4]
  PIN SO[3] 
    ANTENNAPARTIALMETALAREA 23.902 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 115.161 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 1.0088 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 35.0948 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 167.794 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 0.885864 LAYER VIA34 ;
    ANTENNADIFFAREA 0.6 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 11.569 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 56.0317 LAYER METAL4 ;
    ANTENNAGATEAREA 2.6078 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 39.5311 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 189.28 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.972272 LAYER VIA45 ;
  END SO[3]
  PIN SO[2] 
    ANTENNAPARTIALMETALAREA 5.48 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 26.3588 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 94.0459 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 453.566 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.07233 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.25 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3949 LAYER METAL4 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 96.9162 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 469.581 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 29.624 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 142.684 LAYER METAL5 ;
    ANTENNAGATEAREA 0.247 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 216.851 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 1047.25 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA56 ;
  END SO[2]
  PIN SO[1] 
    ANTENNAPARTIALMETALAREA 4.001 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.2448 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.154 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.93314 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 24.203 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 116.609 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.221 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 167.571 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 810.28 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.46443 LAYER VIA56 ;
  END SO[1]
  PIN SO[0] 
    ANTENNAPARTIALMETALAREA 3.005 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.4541 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 56.3881 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 272.431 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAMAXCUTCAR 2.07233 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.25 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.3949 LAYER METAL4 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 59.2583 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 288.446 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 33.76 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 162.578 LAYER METAL5 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 446.859 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 2155.01 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 2.90126 LAYER VIA56 ;
  END SO[0]
  PIN scan_clk 
    ANTENNAPARTIALMETALAREA 0.255 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.22655 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.222 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 1.26022 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 1.534 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.57094 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 1.61865 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 7.93145 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END scan_clk
  PIN scan_rst 
    ANTENNAPARTIALMETALAREA 1.599 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 7.69119 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 2.518 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 12.304 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 7.028 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 33.9971 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1599 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 80.2376 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 389.095 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END scan_rst
  PIN test_mode 
    ANTENNAPARTIALMETALAREA 0.465 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.23665 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.498 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.39778 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0871 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 20.4179 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 101.624 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 1.2434 LAYER VIA34 ;
  END test_mode
  PIN SE 
    ANTENNAPARTIALMETALAREA 0.442 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 2.12602 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 4.181 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 20.303 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1755 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 25.5305 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 124.219 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.617094 LAYER VIA34 ;
  END SE
  PIN RST_N 
    ANTENNAPARTIALMETALAREA 2.041 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 9.81721 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 0.145 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.88985 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 7.356 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 35.5748 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0533 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 192.608 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 933.807 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 2.03189 LAYER VIA45 ;
  END RST_N
  PIN UART_CLK 
    ANTENNAPARTIALMETALAREA 0.241 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 1.15921 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.042 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.20442 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.714 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 3.62674 LAYER METAL4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL4 ; 
    ANTENNAMAXAREACAR 0.654826 LAYER METAL4 ;
    ANTENNAMAXSIDEAREACAR 3.29546 LAYER METAL4 ;
    ANTENNAMAXCUTCAR 0.0353598 LAYER VIA45 ;
  END UART_CLK
  PIN REF_CLK 
    ANTENNAPARTIALMETALAREA 0.141 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 0.67821 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0361 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.384 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 6.84944 LAYER METAL3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 3.0628 LAYER METAL3 ; 
    ANTENNAMAXAREACAR 0.586914 LAYER METAL3 ;
    ANTENNAMAXSIDEAREACAR 2.90598 LAYER METAL3 ;
    ANTENNAMAXCUTCAR 0.0235732 LAYER VIA34 ;
  END REF_CLK
  PIN UART_RX_IN 
    ANTENNAPARTIALMETALAREA 14.706 LAYER METAL2 ;
    ANTENNAPARTIALMETALSIDEAREA 70.7359 LAYER METAL2 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA23 ;
    ANTENNAPARTIALMETALAREA 1.065 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.31505 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 0.35 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.8759 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNAPARTIALMETALAREA 8.468 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 40.9235 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.6617 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 26.6574 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 127.325 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.38746 LAYER VIA56 ;
  END UART_RX_IN
  PIN UART_TX_O 
    ANTENNADIFFAREA 0.524 LAYER METAL3 ; 
    ANTENNAPARTIALMETALAREA 2.342 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.265 LAYER METAL3 ;
  END UART_TX_O
  PIN parity_error 
    ANTENNAPARTIALMETALAREA 3.964 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 19.0668 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNAPARTIALMETALAREA 11.903 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 57.4458 LAYER METAL4 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA45 ;
    ANTENNADIFFAREA 0.6 LAYER METAL5 ; 
    ANTENNAPARTIALMETALAREA 25.114 LAYER METAL5 ;
    ANTENNAPARTIALMETALSIDEAREA 120.991 LAYER METAL5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3185 LAYER METAL5 ; 
    ANTENNAMAXAREACAR 152.779 LAYER METAL5 ;
    ANTENNAMAXSIDEAREACAR 740.156 LAYER METAL5 ;
    ANTENNAMAXCUTCAR 1.80797 LAYER VIA56 ;
  END parity_error
  PIN framing_error 
    ANTENNAPARTIALMETALAREA 2.119 LAYER METAL3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1924 LAYER METAL3 ;
    ANTENNAPARTIALCUTAREA 0.0722 LAYER VIA34 ;
    ANTENNADIFFAREA 0.524 LAYER METAL4 ; 
    ANTENNAPARTIALMETALAREA 7.147 LAYER METAL4 ;
    ANTENNAPARTIALMETALSIDEAREA 34.5695 LAYER METAL4 ;
  END framing_error
END SYS_TOP

END LIBRARY
