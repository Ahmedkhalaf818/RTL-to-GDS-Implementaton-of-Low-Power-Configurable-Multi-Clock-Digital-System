module DLY3X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY4X1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX20M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX18M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX32M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX16M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX40M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX24M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX14M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module TIEHIM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module TIELOM (
	Y, 
	VDD, 
	VSS);
   output Y;
   inout VDD;
   inout VSS;
endmodule

module NAND2X3M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3BX4M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X2M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKAND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X4M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX4M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NAND3X4M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X3M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX8M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKAND2X6M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X4M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XOR2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X8M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND2X6M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MXI2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX8M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR2X3M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X4M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21X6M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND2X4M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X4M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2X8M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI21X8M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X4M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX4M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module CLKNAND2X12M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B2X8M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2X5M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X1M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX2M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module NOR2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB2X8M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI21X4M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MXI2X3M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X4M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI22X4M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI21X3M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX4M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND2X8M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2X4M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module NAND3X6M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND3X6M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX10M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX10M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX2M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module BUFX5M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX8M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKBUFX6M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module DLY1X4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVXLM (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X8M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X6M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module TLATNCAX2M (
	ECK, 
	E, 
	CK, 
	VDD, 
	VSS);
   output ECK;
   input E;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module OR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX2M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX2M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX4M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module INVX4M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module MX4X1M (
	Y, 
	S1, 
	S0, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S1;
   input S0;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO21XLM (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X2M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module XNOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB1X1M (
	Y, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module AOI221XLM (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDHX1M (
	S, 
	CO, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKXOR2X2M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module SDFFRHQX1M (
	SI, 
	SE, 
	RN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NOR3BX4M (
	Y, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module AND3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI31X2M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI222X4M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2BB2XLM (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0N, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0N;
   inout VDD;
   inout VSS;
endmodule

module OAI222X1M (
	Y, 
	C1, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C1;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI211X1M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI32X1M (
	Y, 
	B1, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X1M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI31X1M (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B11X1M (
	Y, 
	C0, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AOI2B1X1M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFHX1M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX14M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX12M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKMX2X2M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module MX2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module ADDFX2M (
	S, 
	CO, 
	CI, 
	B, 
	A, 
	VDD, 
	VSS);
   output S;
   output CO;
   input CI;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AOI21BX2M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module XOR3XLM (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI21BX1M (
	Y, 
	B0N, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0N;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module AND2X1M (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module INVX3M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module AO2B2X2M (
	Y, 
	B1, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module NOR2BX1M (
	Y, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module SDFFRX1M (
	SI, 
	SE, 
	RN, 
	QN, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SI;
   input SE;
   input RN;
   output QN;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module OAI22X1M (
	Y, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module SDFFSQX1M (
	SN, 
	SI, 
	SE, 
	Q, 
	D, 
	CK, 
	VDD, 
	VSS);
   input SN;
   input SI;
   input SE;
   output Q;
   input D;
   input CK;
   inout VDD;
   inout VSS;
endmodule

module NAND4BX1M (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module MXI2X1M (
	Y, 
	S0, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input S0;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module CLKINVX1M (
	Y, 
	A, 
	VDD, 
	VSS);
   output Y;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OR3X1M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X1M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4BXLM (
	Y, 
	D, 
	C, 
	B, 
	AN, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input AN;
   inout VDD;
   inout VSS;
endmodule

module OAI31XLM (
	Y, 
	B0, 
	A2, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A2;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI211X2M (
	Y, 
	C0, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OAI2B1X2M (
	Y, 
	B0, 
	A1N, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1N;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OA21X2M (
	Y, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

module OR3X2M (
	Y, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NOR2XLM (
	Y, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module NAND4X2M (
	Y, 
	D, 
	C, 
	B, 
	A, 
	VDD, 
	VSS);
   output Y;
   input D;
   input C;
   input B;
   input A;
   inout VDD;
   inout VSS;
endmodule

module OAI221X1M (
	Y, 
	C0, 
	B1, 
	B0, 
	A1, 
	A0, 
	VDD, 
	VSS);
   output Y;
   input C0;
   input B1;
   input B0;
   input A1;
   input A0;
   inout VDD;
   inout VSS;
endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : K-2015.06
// Date      : Sat Oct  4 07:24:43 2025
/////////////////////////////////////////////////////////////
module mux2X1_1 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Module instantiations
   MX2X8M U1 (
	.Y(OUT),
	.S0(SEL),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_5 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(SEL),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_4 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN5_scan_rst;
   wire FE_PHN2_scan_rst;
   wire FE_PHN1_RST_N;
   wire FE_PHN0_RST_N;

   // Module instantiations
   DLY4X1M FE_PHC5_scan_rst (
	.Y(FE_PHN5_scan_rst),
	.A(FE_PHN2_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC2_scan_rst (
	.Y(FE_PHN2_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC1_RST_N (
	.Y(FE_PHN1_RST_N),
	.A(FE_PHN0_RST_N), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC0_RST_N (
	.Y(FE_PHN0_RST_N),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U1 (
	.Y(OUT),
	.S0(SEL),
	.B(FE_PHN5_scan_rst),
	.A(FE_PHN1_RST_N), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_3 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(SEL),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_2 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Module instantiations
   MX2X2M U1 (
	.Y(OUT),
	.S0(SEL),
	.B(IN_1),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_0 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN7_scan_rst;
   wire FE_PHN4_scan_rst;

   // Module instantiations
   DLY4X1M FE_PHC7_scan_rst (
	.Y(FE_PHN7_scan_rst),
	.A(FE_PHN4_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC4_scan_rst (
	.Y(FE_PHN4_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X8M U1 (
	.Y(OUT),
	.S0(SEL),
	.B(FE_PHN7_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module mux2X1_6 (
	IN_0, 
	IN_1, 
	SEL, 
	OUT, 
	VDD, 
	VSS);
   input IN_0;
   input IN_1;
   input SEL;
   output OUT;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN6_scan_rst;
   wire FE_PHN3_scan_rst;

   // Module instantiations
   DLY4X1M FE_PHC6_scan_rst (
	.Y(FE_PHN6_scan_rst),
	.A(FE_PHN3_scan_rst), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY4X1M FE_PHC3_scan_rst (
	.Y(FE_PHN3_scan_rst),
	.A(IN_1), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X6M U1 (
	.Y(OUT),
	.S0(SEL),
	.B(FE_PHN6_scan_rst),
	.A(IN_0), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYN_test_0 (
	CLK, 
	RST, 
	SYNC_RST, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output SYNC_RST;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \rst_shift_reg[0] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rst_shift_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\rst_shift_reg[0] ),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \rst_shift_reg_reg[1]  (
	.SI(\rst_shift_reg[0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(\rst_shift_reg[0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RST_SYN_test_1 (
	CLK, 
	RST, 
	SYNC_RST, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   output SYNC_RST;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire \rst_shift_reg[0] ;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \rst_shift_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST),
	.Q(\rst_shift_reg[0] ),
	.D(HTIE_LTIEHI_NET),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M \rst_shift_reg_reg[1]  (
	.SI(\rst_shift_reg[0] ),
	.SE(test_se),
	.RN(RST),
	.Q(SYNC_RST),
	.D(\rst_shift_reg[0] ),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module CLK_gating (
	CLK, 
	CLK_EN, 
	test, 
	Gated_CLK, 
	VDD, 
	VSS);
   input CLK;
   input CLK_EN;
   input test;
   output Gated_CLK;
   inout VDD;
   inout VSS;

   // Internal wires
   wire _2_net_;

   // Module instantiations
   TLATNCAX2M U_LATNCAX2M (
	.ECK(Gated_CLK),
	.E(_2_net_),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U1 (
	.Y(_2_net_),
	.B(test),
	.A(CLK_EN), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module Register_File_test_1 (
	CLK, 
	RST, 
	WrEn, 
	RdEn, 
	Address, 
	WrData, 
	RdData, 
	RdData_valid, 
	REG0, 
	REG1, 
	REG2, 
	REG3, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN0_RST_SYNC_1_mux, 
	CLK_R_M__L5_N4, 
	CLK_R_M__L5_N5, 
	CLK_R_M__L5_N6, 
	CLK_R_M__L5_N7, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input WrEn;
   input RdEn;
   input [3:0] Address;
   input [7:0] WrData;
   output [7:0] RdData;
   output RdData_valid;
   output [7:0] REG0;
   output [7:0] REG1;
   output [7:0] REG2;
   output [7:0] REG3;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN0_RST_SYNC_1_mux;
   input CLK_R_M__L5_N4;
   input CLK_R_M__L5_N5;
   input CLK_R_M__L5_N6;
   input CLK_R_M__L5_N7;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN20_REG1_OP_B_6_;
   wire FE_OFN19_REG0_OP_A_7_;
   wire FE_OFN18_REG0_OP_A_6_;
   wire FE_OFN17_REG0_OP_A_5_;
   wire FE_OFN16_REG0_OP_A_4_;
   wire FE_OFN15_REG0_OP_A_3_;
   wire FE_OFN14_REG0_OP_A_2_;
   wire FE_OFN13_REG1_OP_B_1_;
   wire FE_OFN12_REG1_OP_B_5_;
   wire FE_OFN11_REG1_OP_B_7_;
   wire FE_OFN10_REG1_OP_B_0_;
   wire FE_OFN1_RST_SYNC_1_mux;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire \regfile[15][7] ;
   wire \regfile[15][6] ;
   wire \regfile[15][5] ;
   wire \regfile[15][4] ;
   wire \regfile[15][3] ;
   wire \regfile[15][2] ;
   wire \regfile[15][1] ;
   wire \regfile[15][0] ;
   wire \regfile[14][7] ;
   wire \regfile[14][6] ;
   wire \regfile[14][5] ;
   wire \regfile[14][4] ;
   wire \regfile[14][3] ;
   wire \regfile[14][2] ;
   wire \regfile[14][1] ;
   wire \regfile[14][0] ;
   wire \regfile[13][7] ;
   wire \regfile[13][6] ;
   wire \regfile[13][5] ;
   wire \regfile[13][4] ;
   wire \regfile[13][3] ;
   wire \regfile[13][2] ;
   wire \regfile[13][1] ;
   wire \regfile[13][0] ;
   wire \regfile[12][7] ;
   wire \regfile[12][6] ;
   wire \regfile[12][5] ;
   wire \regfile[12][4] ;
   wire \regfile[12][3] ;
   wire \regfile[12][2] ;
   wire \regfile[12][1] ;
   wire \regfile[12][0] ;
   wire \regfile[11][7] ;
   wire \regfile[11][6] ;
   wire \regfile[11][5] ;
   wire \regfile[11][4] ;
   wire \regfile[11][3] ;
   wire \regfile[11][2] ;
   wire \regfile[11][1] ;
   wire \regfile[11][0] ;
   wire \regfile[10][7] ;
   wire \regfile[10][6] ;
   wire \regfile[10][5] ;
   wire \regfile[10][4] ;
   wire \regfile[10][3] ;
   wire \regfile[10][2] ;
   wire \regfile[10][1] ;
   wire \regfile[10][0] ;
   wire \regfile[9][7] ;
   wire \regfile[9][6] ;
   wire \regfile[9][5] ;
   wire \regfile[9][4] ;
   wire \regfile[9][3] ;
   wire \regfile[9][2] ;
   wire \regfile[9][1] ;
   wire \regfile[9][0] ;
   wire \regfile[8][7] ;
   wire \regfile[8][6] ;
   wire \regfile[8][5] ;
   wire \regfile[8][4] ;
   wire \regfile[8][3] ;
   wire \regfile[8][2] ;
   wire \regfile[8][1] ;
   wire \regfile[8][0] ;
   wire \regfile[7][7] ;
   wire \regfile[7][6] ;
   wire \regfile[7][5] ;
   wire \regfile[7][4] ;
   wire \regfile[7][3] ;
   wire \regfile[7][2] ;
   wire \regfile[7][1] ;
   wire \regfile[7][0] ;
   wire \regfile[6][7] ;
   wire \regfile[6][6] ;
   wire \regfile[6][5] ;
   wire \regfile[6][4] ;
   wire \regfile[6][3] ;
   wire \regfile[6][2] ;
   wire \regfile[6][1] ;
   wire \regfile[6][0] ;
   wire \regfile[5][7] ;
   wire \regfile[5][6] ;
   wire \regfile[5][5] ;
   wire \regfile[5][4] ;
   wire \regfile[5][3] ;
   wire \regfile[5][2] ;
   wire \regfile[5][1] ;
   wire \regfile[5][0] ;
   wire \regfile[4][7] ;
   wire \regfile[4][6] ;
   wire \regfile[4][5] ;
   wire \regfile[4][4] ;
   wire \regfile[4][3] ;
   wire \regfile[4][2] ;
   wire \regfile[4][1] ;
   wire \regfile[4][0] ;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire N43;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n315;
   wire n316;
   wire n317;
   wire n318;
   wire n319;
   wire n320;
   wire n321;
   wire n322;
   wire n323;
   wire n324;
   wire n325;
   wire n326;
   wire n327;
   wire n328;
   wire n329;
   wire n330;
   wire n331;
   wire n332;
   wire n333;
   wire n334;
   wire n336;
   wire n338;
   wire n339;
   wire n340;
   wire n341;
   wire n357;
   wire n358;
   wire n359;
   wire n360;
   wire n361;
   wire n362;
   wire n363;
   wire n364;
   wire n365;
   wire n366;
   wire n371;
   wire n372;
   wire n373;
   wire n374;

   assign N11 = Address[0] ;
   assign N12 = Address[1] ;
   assign N13 = Address[2] ;
   assign N14 = Address[3] ;
   assign test_so2 = \regfile[15][7]  ;
   assign test_so1 = \regfile[12][4]  ;

   // Module instantiations
   BUFX8M FE_OFC20_REG1_OP_B_6_ (
	.Y(REG1[6]),
	.A(FE_OFN20_REG1_OP_B_6_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC19_REG0_OP_A_7_ (
	.Y(REG0[7]),
	.A(FE_OFN19_REG0_OP_A_7_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC18_REG0_OP_A_6_ (
	.Y(REG0[6]),
	.A(FE_OFN18_REG0_OP_A_6_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC17_REG0_OP_A_5_ (
	.Y(REG0[5]),
	.A(FE_OFN17_REG0_OP_A_5_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC16_REG0_OP_A_4_ (
	.Y(REG0[4]),
	.A(FE_OFN16_REG0_OP_A_4_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX10M FE_OFC15_REG0_OP_A_3_ (
	.Y(REG0[3]),
	.A(FE_OFN15_REG0_OP_A_3_), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX2M FE_OFC14_REG0_OP_A_2_ (
	.Y(REG0[2]),
	.A(FE_OFN14_REG0_OP_A_2_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC13_REG1_OP_B_1_ (
	.Y(REG1[1]),
	.A(FE_OFN13_REG1_OP_B_1_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC12_REG1_OP_B_5_ (
	.Y(REG1[5]),
	.A(FE_OFN12_REG1_OP_B_5_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC11_REG1_OP_B_7_ (
	.Y(REG1[7]),
	.A(FE_OFN11_REG1_OP_B_7_), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M FE_OFC10_REG1_OP_B_0_ (
	.Y(REG1[0]),
	.A(FE_OFN10_REG1_OP_B_0_), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKBUFX8M FE_OFC1_RST_SYNC_1_mux (
	.Y(FE_OFN1_RST_SYNC_1_mux),
	.A(RST), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[13][7]  (
	.SI(\regfile[13][6] ),
	.SE(n373),
	.RN(RST),
	.Q(\regfile[13][7] ),
	.D(n298),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[13][6]  (
	.SI(\regfile[13][5] ),
	.SE(n372),
	.RN(RST),
	.Q(\regfile[13][6] ),
	.D(n297),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[13][5]  (
	.SI(\regfile[13][4] ),
	.SE(n371),
	.RN(RST),
	.Q(\regfile[13][5] ),
	.D(n296),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[13][4]  (
	.SI(\regfile[13][3] ),
	.SE(n374),
	.RN(RST),
	.Q(\regfile[13][4] ),
	.D(n295),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[13][3]  (
	.SI(\regfile[13][2] ),
	.SE(n373),
	.RN(RST),
	.Q(\regfile[13][3] ),
	.D(n294),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[13][2]  (
	.SI(\regfile[13][1] ),
	.SE(n372),
	.RN(RST),
	.Q(\regfile[13][2] ),
	.D(n293),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[13][1]  (
	.SI(\regfile[13][0] ),
	.SE(n371),
	.RN(RST),
	.Q(\regfile[13][1] ),
	.D(n292),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[13][0]  (
	.SI(\regfile[12][7] ),
	.SE(n374),
	.RN(RST),
	.Q(\regfile[13][0] ),
	.D(n291),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[9][7]  (
	.SI(\regfile[9][6] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[9][7] ),
	.D(n266),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[9][6]  (
	.SI(\regfile[9][5] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[9][6] ),
	.D(n265),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[9][5]  (
	.SI(\regfile[9][4] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[9][5] ),
	.D(n264),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[9][4]  (
	.SI(\regfile[9][3] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[9][4] ),
	.D(n263),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[9][3]  (
	.SI(\regfile[9][2] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[9][3] ),
	.D(n262),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[9][2]  (
	.SI(\regfile[9][1] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[9][2] ),
	.D(n261),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[9][1]  (
	.SI(\regfile[9][0] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[9][1] ),
	.D(n260),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[9][0]  (
	.SI(\regfile[8][7] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[9][0] ),
	.D(n259),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[5][7]  (
	.SI(\regfile[5][6] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[5][7] ),
	.D(n234),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[5][6]  (
	.SI(\regfile[5][5] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[5][6] ),
	.D(n233),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[5][5]  (
	.SI(\regfile[5][4] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[5][5] ),
	.D(n232),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[5][4]  (
	.SI(\regfile[5][3] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[5][4] ),
	.D(n231),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[5][3]  (
	.SI(\regfile[5][2] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[5][3] ),
	.D(n230),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[5][2]  (
	.SI(\regfile[5][1] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[5][2] ),
	.D(n229),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[5][1]  (
	.SI(\regfile[5][0] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[5][1] ),
	.D(n228),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[5][0]  (
	.SI(\regfile[4][7] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[5][0] ),
	.D(n227),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[15][7]  (
	.SI(\regfile[15][6] ),
	.SE(n373),
	.RN(RST),
	.Q(\regfile[15][7] ),
	.D(n314),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[15][6]  (
	.SI(\regfile[15][5] ),
	.SE(n372),
	.RN(RST),
	.Q(\regfile[15][6] ),
	.D(n313),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[15][5]  (
	.SI(\regfile[15][4] ),
	.SE(n371),
	.RN(RST),
	.Q(\regfile[15][5] ),
	.D(n312),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[15][4]  (
	.SI(\regfile[15][3] ),
	.SE(n374),
	.RN(RST),
	.Q(\regfile[15][4] ),
	.D(n311),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[15][3]  (
	.SI(\regfile[15][2] ),
	.SE(n373),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(\regfile[15][3] ),
	.D(n310),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[15][2]  (
	.SI(\regfile[15][1] ),
	.SE(n372),
	.RN(RST),
	.Q(\regfile[15][2] ),
	.D(n309),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[15][1]  (
	.SI(\regfile[15][0] ),
	.SE(n371),
	.RN(RST),
	.Q(\regfile[15][1] ),
	.D(n308),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[15][0]  (
	.SI(\regfile[14][7] ),
	.SE(n374),
	.RN(RST),
	.Q(\regfile[15][0] ),
	.D(n307),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[11][7]  (
	.SI(\regfile[11][6] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[11][7] ),
	.D(n282),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[11][6]  (
	.SI(\regfile[11][5] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[11][6] ),
	.D(n281),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[11][5]  (
	.SI(\regfile[11][4] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[11][5] ),
	.D(n280),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[11][4]  (
	.SI(\regfile[11][3] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[11][4] ),
	.D(n279),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[11][3]  (
	.SI(\regfile[11][2] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[11][3] ),
	.D(n278),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[11][2]  (
	.SI(\regfile[11][1] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[11][2] ),
	.D(n277),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[11][1]  (
	.SI(\regfile[11][0] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[11][1] ),
	.D(n276),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[11][0]  (
	.SI(\regfile[10][7] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[11][0] ),
	.D(n275),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[7][7]  (
	.SI(\regfile[7][6] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[7][7] ),
	.D(n250),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[7][6]  (
	.SI(\regfile[7][5] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[7][6] ),
	.D(n249),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[7][5]  (
	.SI(\regfile[7][4] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[7][5] ),
	.D(n248),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[7][4]  (
	.SI(\regfile[7][3] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[7][4] ),
	.D(n247),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[7][3]  (
	.SI(\regfile[7][2] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[7][3] ),
	.D(n246),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[7][2]  (
	.SI(\regfile[7][1] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[7][2] ),
	.D(n245),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[7][1]  (
	.SI(\regfile[7][0] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[7][1] ),
	.D(n244),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[7][0]  (
	.SI(\regfile[6][7] ),
	.SE(n374),
	.RN(RST),
	.Q(\regfile[7][0] ),
	.D(n243),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[14][7]  (
	.SI(\regfile[14][6] ),
	.SE(n373),
	.RN(RST),
	.Q(\regfile[14][7] ),
	.D(n306),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[14][6]  (
	.SI(\regfile[14][5] ),
	.SE(n372),
	.RN(RST),
	.Q(\regfile[14][6] ),
	.D(n305),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[14][5]  (
	.SI(\regfile[14][4] ),
	.SE(n371),
	.RN(RST),
	.Q(\regfile[14][5] ),
	.D(n304),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[14][4]  (
	.SI(\regfile[14][3] ),
	.SE(n374),
	.RN(RST),
	.Q(\regfile[14][4] ),
	.D(n303),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[14][3]  (
	.SI(\regfile[14][2] ),
	.SE(n373),
	.RN(RST),
	.Q(\regfile[14][3] ),
	.D(n302),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[14][2]  (
	.SI(\regfile[14][1] ),
	.SE(n372),
	.RN(RST),
	.Q(\regfile[14][2] ),
	.D(n301),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[14][1]  (
	.SI(\regfile[14][0] ),
	.SE(n371),
	.RN(RST),
	.Q(\regfile[14][1] ),
	.D(n300),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[14][0]  (
	.SI(\regfile[13][7] ),
	.SE(n374),
	.RN(RST),
	.Q(\regfile[14][0] ),
	.D(n299),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[10][7]  (
	.SI(\regfile[10][6] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[10][7] ),
	.D(n274),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[10][6]  (
	.SI(\regfile[10][5] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[10][6] ),
	.D(n273),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[10][5]  (
	.SI(\regfile[10][4] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[10][5] ),
	.D(n272),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[10][4]  (
	.SI(\regfile[10][3] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[10][4] ),
	.D(n271),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[10][3]  (
	.SI(\regfile[10][2] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[10][3] ),
	.D(n270),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[10][2]  (
	.SI(\regfile[10][1] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[10][2] ),
	.D(n269),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[10][1]  (
	.SI(\regfile[10][0] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[10][1] ),
	.D(n268),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[10][0]  (
	.SI(\regfile[9][7] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[10][0] ),
	.D(n267),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[6][7]  (
	.SI(\regfile[6][6] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[6][7] ),
	.D(n242),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[6][6]  (
	.SI(\regfile[6][5] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[6][6] ),
	.D(n241),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[6][5]  (
	.SI(\regfile[6][4] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[6][5] ),
	.D(n240),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[6][4]  (
	.SI(\regfile[6][3] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[6][4] ),
	.D(n239),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[6][3]  (
	.SI(\regfile[6][2] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[6][3] ),
	.D(n238),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[6][2]  (
	.SI(\regfile[6][1] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[6][2] ),
	.D(n237),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[6][1]  (
	.SI(\regfile[6][0] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[6][1] ),
	.D(n236),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[6][0]  (
	.SI(\regfile[5][7] ),
	.SE(n374),
	.RN(RST),
	.Q(\regfile[6][0] ),
	.D(n235),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[12][7]  (
	.SI(\regfile[12][6] ),
	.SE(n373),
	.RN(RST),
	.Q(\regfile[12][7] ),
	.D(n290),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[12][6]  (
	.SI(\regfile[12][5] ),
	.SE(n372),
	.RN(RST),
	.Q(\regfile[12][6] ),
	.D(n289),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[12][5]  (
	.SI(test_si3),
	.SE(n371),
	.RN(RST),
	.Q(\regfile[12][5] ),
	.D(n288),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \regfile_reg[12][4]  (
	.SI(\regfile[12][3] ),
	.SE(n374),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(\regfile[12][4] ),
	.D(n287),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[12][3]  (
	.SI(\regfile[12][2] ),
	.SE(n373),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(\regfile[12][3] ),
	.D(n286),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[12][2]  (
	.SI(\regfile[12][1] ),
	.SE(n372),
	.RN(RST),
	.Q(\regfile[12][2] ),
	.D(n285),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[12][1]  (
	.SI(\regfile[12][0] ),
	.SE(n371),
	.RN(RST),
	.Q(\regfile[12][1] ),
	.D(n284),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[12][0]  (
	.SI(\regfile[11][7] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[12][0] ),
	.D(n283),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[8][7]  (
	.SI(\regfile[8][6] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[8][7] ),
	.D(n258),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[8][6]  (
	.SI(\regfile[8][5] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[8][6] ),
	.D(n257),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[8][5]  (
	.SI(\regfile[8][4] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[8][5] ),
	.D(n256),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[8][4]  (
	.SI(\regfile[8][3] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[8][4] ),
	.D(n255),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[8][3]  (
	.SI(\regfile[8][2] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[8][3] ),
	.D(n254),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[8][2]  (
	.SI(\regfile[8][1] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[8][2] ),
	.D(n253),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[8][1]  (
	.SI(\regfile[8][0] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[8][1] ),
	.D(n252),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[8][0]  (
	.SI(\regfile[7][7] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[8][0] ),
	.D(n251),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[4][7]  (
	.SI(\regfile[4][6] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[4][7] ),
	.D(n226),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[4][6]  (
	.SI(\regfile[4][5] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[4][6] ),
	.D(n225),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[4][5]  (
	.SI(\regfile[4][4] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[4][5] ),
	.D(n224),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[4][4]  (
	.SI(\regfile[4][3] ),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[4][4] ),
	.D(n223),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[4][3]  (
	.SI(\regfile[4][2] ),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[4][3] ),
	.D(n222),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[4][2]  (
	.SI(\regfile[4][1] ),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[4][2] ),
	.D(n221),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[4][1]  (
	.SI(\regfile[4][0] ),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[4][1] ),
	.D(n220),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[4][0]  (
	.SI(REG3[7]),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(\regfile[4][0] ),
	.D(n219),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[7]  (
	.SI(RdData[6]),
	.SE(n373),
	.RN(RST),
	.Q(RdData[7]),
	.D(n186),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[6]  (
	.SI(RdData[5]),
	.SE(n372),
	.RN(RST),
	.Q(RdData[6]),
	.D(n185),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[5]  (
	.SI(RdData[4]),
	.SE(n371),
	.RN(RST),
	.Q(RdData[5]),
	.D(n184),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[4]  (
	.SI(RdData[3]),
	.SE(n374),
	.RN(RST),
	.Q(RdData[4]),
	.D(n183),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[3]  (
	.SI(RdData[2]),
	.SE(n373),
	.RN(RST),
	.Q(RdData[3]),
	.D(n182),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[2]  (
	.SI(RdData[1]),
	.SE(n372),
	.RN(RST),
	.Q(RdData[2]),
	.D(n181),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[1]  (
	.SI(RdData[0]),
	.SE(n371),
	.RN(RST),
	.Q(RdData[1]),
	.D(n180),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RdData_reg[0]  (
	.SI(test_si1),
	.SE(n374),
	.RN(RST),
	.Q(RdData[0]),
	.D(n179),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \regfile_reg[1][6]  (
	.SI(REG1[5]),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(FE_OFN20_REG1_OP_B_6_),
	.D(n201),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \regfile_reg[0][7]  (
	.SI(REG0[6]),
	.SE(n372),
	.RN(RST),
	.Q(FE_OFN19_REG0_OP_A_7_),
	.D(n194),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \regfile_reg[0][6]  (
	.SI(REG0[5]),
	.SE(n371),
	.RN(RST),
	.Q(FE_OFN18_REG0_OP_A_6_),
	.D(n193),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \regfile_reg[0][5]  (
	.SI(REG0[4]),
	.SE(n374),
	.RN(RST),
	.Q(FE_OFN17_REG0_OP_A_5_),
	.D(n192),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \regfile_reg[0][4]  (
	.SI(REG0[3]),
	.SE(n373),
	.RN(RST),
	.Q(FE_OFN16_REG0_OP_A_4_),
	.D(n191),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \regfile_reg[0][3]  (
	.SI(REG0[2]),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(FE_OFN15_REG0_OP_A_3_),
	.D(n190),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[0][2]  (
	.SI(REG0[1]),
	.SE(n371),
	.RN(RST),
	.Q(FE_OFN14_REG0_OP_A_2_),
	.D(n189),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[0][1]  (
	.SI(REG0[0]),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(REG0[1]),
	.D(n188),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[0][0]  (
	.SI(RdData_valid),
	.SE(n373),
	.RN(RST),
	.Q(REG0[0]),
	.D(n187),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[2][1]  (
	.SI(REG2[0]),
	.SE(n372),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(REG2[1]),
	.D(n204),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[3][0]  (
	.SI(REG2[7]),
	.SE(n371),
	.RN(RST),
	.Q(REG3[0]),
	.D(n211),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \regfile_reg[2][0]  (
	.SN(RST),
	.SI(REG1[7]),
	.SE(test_se),
	.Q(REG2[0]),
	.D(n203),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \regfile_reg[1][1]  (
	.SI(REG1[0]),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(FE_OFN13_REG1_OP_B_1_),
	.D(n196),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \regfile_reg[1][5]  (
	.SI(REG1[4]),
	.SE(n373),
	.RN(RST),
	.Q(FE_OFN12_REG1_OP_B_5_),
	.D(n200),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \regfile_reg[1][4]  (
	.SI(REG1[3]),
	.SE(n372),
	.RN(RST),
	.Q(REG1[4]),
	.D(n199),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX2M \regfile_reg[1][7]  (
	.SI(REG1[6]),
	.SE(n371),
	.RN(RST),
	.Q(FE_OFN11_REG1_OP_B_7_),
	.D(n202),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \regfile_reg[1][3]  (
	.SI(REG1[2]),
	.SE(n374),
	.RN(RST),
	.Q(REG1[3]),
	.D(n198),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \regfile_reg[1][2]  (
	.SI(REG1[1]),
	.SE(n373),
	.RN(RST),
	.Q(REG1[2]),
	.D(n197),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX4M \regfile_reg[1][0]  (
	.SI(REG0[7]),
	.SE(n372),
	.RN(RST),
	.Q(FE_OFN10_REG1_OP_B_0_),
	.D(n195),
	.CK(CLK_R_M__L5_N6), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M RdData_valid_reg (
	.SI(RdData[7]),
	.SE(n371),
	.RN(RST),
	.Q(RdData_valid),
	.D(n178),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \regfile_reg[3][5]  (
	.SN(RST),
	.SI(REG3[4]),
	.SE(n371),
	.Q(REG3[5]),
	.D(n216),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[3][7]  (
	.SI(REG3[6]),
	.SE(n374),
	.RN(RST),
	.Q(REG3[7]),
	.D(n218),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[3][4]  (
	.SI(REG3[3]),
	.SE(n373),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(REG3[4]),
	.D(n215),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[3][6]  (
	.SI(REG3[5]),
	.SE(n372),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(REG3[6]),
	.D(n217),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[3][3]  (
	.SI(REG3[2]),
	.SE(n371),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(REG3[3]),
	.D(n214),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[3][2]  (
	.SI(REG3[1]),
	.SE(n374),
	.RN(FE_OFN1_RST_SYNC_1_mux),
	.Q(REG3[2]),
	.D(n213),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[3][1]  (
	.SI(REG3[0]),
	.SE(n373),
	.RN(RST),
	.Q(REG3[1]),
	.D(n212),
	.CK(CLK_R_M__L5_N7), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[2][2]  (
	.SI(REG2[1]),
	.SE(n372),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(REG2[2]),
	.D(n205),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \regfile_reg[2][7]  (
	.SN(RST),
	.SI(REG2[6]),
	.SE(n374),
	.Q(REG2[7]),
	.D(n210),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[2][6]  (
	.SI(REG2[5]),
	.SE(n371),
	.RN(RST),
	.Q(REG2[6]),
	.D(n209),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[2][5]  (
	.SI(REG2[4]),
	.SE(n374),
	.RN(RST),
	.Q(REG2[5]),
	.D(n208),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[2][4]  (
	.SI(REG2[3]),
	.SE(n373),
	.RN(RST),
	.Q(REG2[4]),
	.D(n207),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \regfile_reg[2][3]  (
	.SI(test_si2),
	.SE(n372),
	.RN(RST),
	.Q(REG2[3]),
	.D(n206),
	.CK(CLK_R_M__L5_N5), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U140 (
	.Y(n365),
	.A(WrData[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U141 (
	.Y(n366),
	.A(WrData[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U142 (
	.Y(n158),
	.B(N13),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U143 (
	.Y(n153),
	.B(N13),
	.A(n336), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U144 (
	.Y(n338),
	.A(n340), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U145 (
	.Y(n336),
	.A(n341), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U146 (
	.Y(n339),
	.A(n340), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U149 (
	.Y(n362),
	.A(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U150 (
	.Y(n357),
	.A(WrData[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U151 (
	.Y(n361),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U162 (
	.Y(n155),
	.B(n153),
	.A(n156), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U163 (
	.Y(n157),
	.B(n154),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U164 (
	.Y(n159),
	.B(n156),
	.A(n158), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U165 (
	.Y(n160),
	.B(n154),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U166 (
	.Y(n162),
	.B(n156),
	.A(n161), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U167 (
	.Y(n163),
	.B(n154),
	.A(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U168 (
	.Y(n166),
	.B(n156),
	.A(n164), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U169 (
	.Y(n167),
	.B(n153),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U170 (
	.Y(n169),
	.B(n153),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U171 (
	.Y(n171),
	.B(n158),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U172 (
	.Y(n172),
	.B(n158),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U173 (
	.Y(n173),
	.B(n161),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U174 (
	.Y(n174),
	.B(n161),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U175 (
	.Y(n175),
	.B(n164),
	.A(n168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U176 (
	.Y(n177),
	.B(n164),
	.A(n170), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U177 (
	.Y(n152),
	.B(n154),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U178 (
	.Y(n151),
	.B(n362),
	.A(RdEn), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U179 (
	.Y(n150),
	.B(RdEn),
	.A(n362), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U180 (
	.Y(n154),
	.B(n340),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U181 (
	.Y(n156),
	.B(N11),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U182 (
	.Y(n168),
	.B(n340),
	.A(n176), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U183 (
	.Y(n170),
	.B(N11),
	.A(n176), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U184 (
	.Y(n358),
	.A(WrData[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U185 (
	.Y(n359),
	.A(WrData[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U186 (
	.Y(n360),
	.A(WrData[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U187 (
	.Y(n364),
	.A(WrData[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U188 (
	.Y(n363),
	.A(WrData[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U194 (
	.Y(n187),
	.B1(n357),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U195 (
	.Y(n188),
	.B1(n358),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U196 (
	.Y(n189),
	.B1(n359),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U197 (
	.Y(n190),
	.B1(n360),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U198 (
	.Y(n191),
	.B1(n364),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U199 (
	.Y(n192),
	.B1(n365),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U200 (
	.Y(n193),
	.B1(n363),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U201 (
	.Y(n194),
	.B1(n366),
	.B0(n152),
	.A1N(n152),
	.A0N(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U202 (
	.Y(n204),
	.B1(n157),
	.B0(n358),
	.A1N(n157),
	.A0N(REG2[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U203 (
	.Y(n205),
	.B1(n157),
	.B0(n359),
	.A1N(n157),
	.A0N(REG2[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U204 (
	.Y(n206),
	.B1(n157),
	.B0(n360),
	.A1N(n157),
	.A0N(REG2[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U205 (
	.Y(n207),
	.B1(n157),
	.B0(n364),
	.A1N(n157),
	.A0N(REG2[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U206 (
	.Y(n208),
	.B1(n157),
	.B0(n365),
	.A1N(n157),
	.A0N(REG2[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U207 (
	.Y(n209),
	.B1(n157),
	.B0(n363),
	.A1N(n157),
	.A0N(REG2[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U208 (
	.Y(n211),
	.B1(n159),
	.B0(n357),
	.A1N(n159),
	.A0N(REG3[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U209 (
	.Y(n212),
	.B1(n159),
	.B0(n358),
	.A1N(n159),
	.A0N(REG3[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U210 (
	.Y(n213),
	.B1(n159),
	.B0(n359),
	.A1N(n159),
	.A0N(REG3[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U211 (
	.Y(n214),
	.B1(n159),
	.B0(n360),
	.A1N(n159),
	.A0N(REG3[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U212 (
	.Y(n215),
	.B1(n159),
	.B0(n364),
	.A1N(n159),
	.A0N(REG3[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U213 (
	.Y(n217),
	.B1(n159),
	.B0(n363),
	.A1N(n159),
	.A0N(REG3[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U214 (
	.Y(n218),
	.B1(n159),
	.B0(n366),
	.A1N(n159),
	.A0N(REG3[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U215 (
	.Y(n195),
	.B1(n155),
	.B0(n357),
	.A1N(n155),
	.A0N(REG1[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U216 (
	.Y(n196),
	.B1(n155),
	.B0(n358),
	.A1N(n155),
	.A0N(REG1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U217 (
	.Y(n197),
	.B1(n155),
	.B0(n359),
	.A1N(n155),
	.A0N(REG1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U218 (
	.Y(n198),
	.B1(n155),
	.B0(n360),
	.A1N(n155),
	.A0N(REG1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U219 (
	.Y(n199),
	.B1(n155),
	.B0(n364),
	.A1N(n155),
	.A0N(REG1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U220 (
	.Y(n200),
	.B1(n155),
	.B0(n365),
	.A1N(n155),
	.A0N(REG1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U221 (
	.Y(n201),
	.B1(n155),
	.B0(n363),
	.A1N(n155),
	.A0N(REG1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U222 (
	.Y(n202),
	.B1(n155),
	.B0(n366),
	.A1N(n155),
	.A0N(REG1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U223 (
	.Y(n251),
	.B1(n167),
	.B0(n357),
	.A1N(n167),
	.A0N(\regfile[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U224 (
	.Y(n252),
	.B1(n167),
	.B0(n358),
	.A1N(n167),
	.A0N(\regfile[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U225 (
	.Y(n253),
	.B1(n167),
	.B0(n359),
	.A1N(n167),
	.A0N(\regfile[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U226 (
	.Y(n254),
	.B1(n167),
	.B0(n360),
	.A1N(n167),
	.A0N(\regfile[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U227 (
	.Y(n255),
	.B1(n167),
	.B0(n364),
	.A1N(n167),
	.A0N(\regfile[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U228 (
	.Y(n256),
	.B1(n167),
	.B0(n365),
	.A1N(n167),
	.A0N(\regfile[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U229 (
	.Y(n257),
	.B1(n167),
	.B0(n363),
	.A1N(n167),
	.A0N(\regfile[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U230 (
	.Y(n258),
	.B1(n167),
	.B0(n366),
	.A1N(n167),
	.A0N(\regfile[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U231 (
	.Y(n259),
	.B1(n169),
	.B0(n357),
	.A1N(n169),
	.A0N(\regfile[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U232 (
	.Y(n260),
	.B1(n169),
	.B0(n358),
	.A1N(n169),
	.A0N(\regfile[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U233 (
	.Y(n261),
	.B1(n169),
	.B0(n359),
	.A1N(n169),
	.A0N(\regfile[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U234 (
	.Y(n262),
	.B1(n169),
	.B0(n360),
	.A1N(n169),
	.A0N(\regfile[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U235 (
	.Y(n263),
	.B1(n169),
	.B0(n364),
	.A1N(n169),
	.A0N(\regfile[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U236 (
	.Y(n264),
	.B1(n169),
	.B0(n365),
	.A1N(n169),
	.A0N(\regfile[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U237 (
	.Y(n265),
	.B1(n169),
	.B0(n363),
	.A1N(n169),
	.A0N(\regfile[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U238 (
	.Y(n266),
	.B1(n169),
	.B0(n366),
	.A1N(n169),
	.A0N(\regfile[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U239 (
	.Y(n267),
	.B1(n171),
	.B0(n357),
	.A1N(n171),
	.A0N(\regfile[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U240 (
	.Y(n268),
	.B1(n171),
	.B0(n358),
	.A1N(n171),
	.A0N(\regfile[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U241 (
	.Y(n269),
	.B1(n171),
	.B0(n359),
	.A1N(n171),
	.A0N(\regfile[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U242 (
	.Y(n270),
	.B1(n171),
	.B0(n360),
	.A1N(n171),
	.A0N(\regfile[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U243 (
	.Y(n271),
	.B1(n171),
	.B0(n364),
	.A1N(n171),
	.A0N(\regfile[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U244 (
	.Y(n272),
	.B1(n171),
	.B0(n365),
	.A1N(n171),
	.A0N(\regfile[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U245 (
	.Y(n273),
	.B1(n171),
	.B0(n363),
	.A1N(n171),
	.A0N(\regfile[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U246 (
	.Y(n274),
	.B1(n171),
	.B0(n366),
	.A1N(n171),
	.A0N(\regfile[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U247 (
	.Y(n275),
	.B1(n172),
	.B0(n357),
	.A1N(n172),
	.A0N(\regfile[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U248 (
	.Y(n276),
	.B1(n172),
	.B0(n358),
	.A1N(n172),
	.A0N(\regfile[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U249 (
	.Y(n277),
	.B1(n172),
	.B0(n359),
	.A1N(n172),
	.A0N(\regfile[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U250 (
	.Y(n278),
	.B1(n172),
	.B0(n360),
	.A1N(n172),
	.A0N(\regfile[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U251 (
	.Y(n279),
	.B1(n172),
	.B0(n364),
	.A1N(n172),
	.A0N(\regfile[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U252 (
	.Y(n280),
	.B1(n172),
	.B0(n365),
	.A1N(n172),
	.A0N(\regfile[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U253 (
	.Y(n281),
	.B1(n172),
	.B0(n363),
	.A1N(n172),
	.A0N(\regfile[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U254 (
	.Y(n282),
	.B1(n172),
	.B0(n366),
	.A1N(n172),
	.A0N(\regfile[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U255 (
	.Y(n203),
	.B1(n157),
	.B0(n357),
	.A1N(n157),
	.A0N(REG2[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U256 (
	.Y(n210),
	.B1(n157),
	.B0(n366),
	.A1N(n157),
	.A0N(REG2[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U257 (
	.Y(n216),
	.B1(n159),
	.B0(n365),
	.A1N(n159),
	.A0N(REG3[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U258 (
	.Y(n219),
	.B1(n160),
	.B0(n357),
	.A1N(n160),
	.A0N(\regfile[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U259 (
	.Y(n220),
	.B1(n160),
	.B0(n358),
	.A1N(n160),
	.A0N(\regfile[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U260 (
	.Y(n221),
	.B1(n160),
	.B0(n359),
	.A1N(n160),
	.A0N(\regfile[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U261 (
	.Y(n222),
	.B1(n160),
	.B0(n360),
	.A1N(n160),
	.A0N(\regfile[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U262 (
	.Y(n223),
	.B1(n160),
	.B0(n364),
	.A1N(n160),
	.A0N(\regfile[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U263 (
	.Y(n224),
	.B1(n160),
	.B0(n365),
	.A1N(n160),
	.A0N(\regfile[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U264 (
	.Y(n225),
	.B1(n160),
	.B0(n363),
	.A1N(n160),
	.A0N(\regfile[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U265 (
	.Y(n226),
	.B1(n160),
	.B0(n366),
	.A1N(n160),
	.A0N(\regfile[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U266 (
	.Y(n227),
	.B1(n162),
	.B0(n357),
	.A1N(n162),
	.A0N(\regfile[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U267 (
	.Y(n228),
	.B1(n162),
	.B0(n358),
	.A1N(n162),
	.A0N(\regfile[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U268 (
	.Y(n229),
	.B1(n162),
	.B0(n359),
	.A1N(n162),
	.A0N(\regfile[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U269 (
	.Y(n230),
	.B1(n162),
	.B0(n360),
	.A1N(n162),
	.A0N(\regfile[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U270 (
	.Y(n231),
	.B1(n162),
	.B0(n364),
	.A1N(n162),
	.A0N(\regfile[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U271 (
	.Y(n232),
	.B1(n162),
	.B0(n365),
	.A1N(n162),
	.A0N(\regfile[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U272 (
	.Y(n233),
	.B1(n162),
	.B0(n363),
	.A1N(n162),
	.A0N(\regfile[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U273 (
	.Y(n234),
	.B1(n162),
	.B0(n366),
	.A1N(n162),
	.A0N(\regfile[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U274 (
	.Y(n235),
	.B1(n163),
	.B0(n357),
	.A1N(n163),
	.A0N(\regfile[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U275 (
	.Y(n236),
	.B1(n163),
	.B0(n358),
	.A1N(n163),
	.A0N(\regfile[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U276 (
	.Y(n237),
	.B1(n163),
	.B0(n359),
	.A1N(n163),
	.A0N(\regfile[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U277 (
	.Y(n238),
	.B1(n163),
	.B0(n360),
	.A1N(n163),
	.A0N(\regfile[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U278 (
	.Y(n239),
	.B1(n163),
	.B0(n364),
	.A1N(n163),
	.A0N(\regfile[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U279 (
	.Y(n240),
	.B1(n163),
	.B0(n365),
	.A1N(n163),
	.A0N(\regfile[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U280 (
	.Y(n241),
	.B1(n163),
	.B0(n363),
	.A1N(n163),
	.A0N(\regfile[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U281 (
	.Y(n242),
	.B1(n163),
	.B0(n366),
	.A1N(n163),
	.A0N(\regfile[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U282 (
	.Y(n243),
	.B1(n166),
	.B0(n357),
	.A1N(n166),
	.A0N(\regfile[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U283 (
	.Y(n244),
	.B1(n166),
	.B0(n358),
	.A1N(n166),
	.A0N(\regfile[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U284 (
	.Y(n245),
	.B1(n166),
	.B0(n359),
	.A1N(n166),
	.A0N(\regfile[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U285 (
	.Y(n246),
	.B1(n166),
	.B0(n360),
	.A1N(n166),
	.A0N(\regfile[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U286 (
	.Y(n247),
	.B1(n166),
	.B0(n364),
	.A1N(n166),
	.A0N(\regfile[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U287 (
	.Y(n248),
	.B1(n166),
	.B0(n365),
	.A1N(n166),
	.A0N(\regfile[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U288 (
	.Y(n249),
	.B1(n166),
	.B0(n363),
	.A1N(n166),
	.A0N(\regfile[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U289 (
	.Y(n250),
	.B1(n166),
	.B0(n366),
	.A1N(n166),
	.A0N(\regfile[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U290 (
	.Y(n283),
	.B1(n173),
	.B0(n357),
	.A1N(n173),
	.A0N(\regfile[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U291 (
	.Y(n284),
	.B1(n173),
	.B0(n358),
	.A1N(n173),
	.A0N(\regfile[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U292 (
	.Y(n285),
	.B1(n173),
	.B0(n359),
	.A1N(n173),
	.A0N(\regfile[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U293 (
	.Y(n286),
	.B1(n173),
	.B0(n360),
	.A1N(n173),
	.A0N(\regfile[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U294 (
	.Y(n287),
	.B1(n173),
	.B0(n364),
	.A1N(n173),
	.A0N(\regfile[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U295 (
	.Y(n288),
	.B1(n173),
	.B0(n365),
	.A1N(n173),
	.A0N(\regfile[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U296 (
	.Y(n289),
	.B1(n173),
	.B0(n363),
	.A1N(n173),
	.A0N(\regfile[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U297 (
	.Y(n290),
	.B1(n173),
	.B0(n366),
	.A1N(n173),
	.A0N(\regfile[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U298 (
	.Y(n291),
	.B1(n174),
	.B0(n357),
	.A1N(n174),
	.A0N(\regfile[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U299 (
	.Y(n292),
	.B1(n174),
	.B0(n358),
	.A1N(n174),
	.A0N(\regfile[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U300 (
	.Y(n293),
	.B1(n174),
	.B0(n359),
	.A1N(n174),
	.A0N(\regfile[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U301 (
	.Y(n294),
	.B1(n174),
	.B0(n360),
	.A1N(n174),
	.A0N(\regfile[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U302 (
	.Y(n295),
	.B1(n174),
	.B0(n364),
	.A1N(n174),
	.A0N(\regfile[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U303 (
	.Y(n296),
	.B1(n174),
	.B0(n365),
	.A1N(n174),
	.A0N(\regfile[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U304 (
	.Y(n297),
	.B1(n174),
	.B0(n363),
	.A1N(n174),
	.A0N(\regfile[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U305 (
	.Y(n298),
	.B1(n174),
	.B0(n366),
	.A1N(n174),
	.A0N(\regfile[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U306 (
	.Y(n299),
	.B1(n175),
	.B0(n357),
	.A1N(n175),
	.A0N(\regfile[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U307 (
	.Y(n300),
	.B1(n175),
	.B0(n358),
	.A1N(n175),
	.A0N(\regfile[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U308 (
	.Y(n301),
	.B1(n175),
	.B0(n359),
	.A1N(n175),
	.A0N(\regfile[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U309 (
	.Y(n302),
	.B1(n175),
	.B0(n360),
	.A1N(n175),
	.A0N(\regfile[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U310 (
	.Y(n303),
	.B1(n175),
	.B0(n364),
	.A1N(n175),
	.A0N(\regfile[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U311 (
	.Y(n304),
	.B1(n175),
	.B0(n365),
	.A1N(n175),
	.A0N(\regfile[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U312 (
	.Y(n305),
	.B1(n175),
	.B0(n363),
	.A1N(n175),
	.A0N(\regfile[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U313 (
	.Y(n306),
	.B1(n175),
	.B0(n366),
	.A1N(n175),
	.A0N(\regfile[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U314 (
	.Y(n307),
	.B1(n177),
	.B0(n357),
	.A1N(n177),
	.A0N(\regfile[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U315 (
	.Y(n308),
	.B1(n177),
	.B0(n358),
	.A1N(n177),
	.A0N(\regfile[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U316 (
	.Y(n309),
	.B1(n177),
	.B0(n359),
	.A1N(n177),
	.A0N(\regfile[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U317 (
	.Y(n310),
	.B1(n177),
	.B0(n360),
	.A1N(n177),
	.A0N(\regfile[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U318 (
	.Y(n311),
	.B1(n177),
	.B0(n364),
	.A1N(n177),
	.A0N(\regfile[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U319 (
	.Y(n312),
	.B1(n177),
	.B0(n365),
	.A1N(n177),
	.A0N(\regfile[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U320 (
	.Y(n313),
	.B1(n177),
	.B0(n363),
	.A1N(n177),
	.A0N(\regfile[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U321 (
	.Y(n314),
	.B1(n177),
	.B0(n366),
	.A1N(n177),
	.A0N(\regfile[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U322 (
	.Y(n165),
	.B(N14),
	.AN(n150), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U323 (
	.Y(n176),
	.B(n150),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U324 (
	.Y(n179),
	.B1(n151),
	.B0(RdData[0]),
	.A1(n361),
	.A0(N43), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U325 (
	.Y(N43),
	.S1(N13),
	.S0(N14),
	.D(n138),
	.C(n140),
	.B(n139),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U326 (
	.Y(n141),
	.S1(n336),
	.S0(N11),
	.D(REG3[0]),
	.C(REG2[0]),
	.B(REG1[0]),
	.A(REG0[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U327 (
	.Y(n139),
	.S1(n336),
	.S0(N11),
	.D(\regfile[11][0] ),
	.C(\regfile[10][0] ),
	.B(\regfile[9][0] ),
	.A(\regfile[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U328 (
	.Y(n180),
	.B1(n151),
	.B0(RdData[1]),
	.A1(n361),
	.A0(N42), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U329 (
	.Y(N42),
	.S1(N13),
	.S0(N14),
	.D(n142),
	.C(n144),
	.B(n143),
	.A(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U330 (
	.Y(n143),
	.S1(n336),
	.S0(N11),
	.D(\regfile[11][1] ),
	.C(\regfile[10][1] ),
	.B(\regfile[9][1] ),
	.A(\regfile[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U331 (
	.Y(n142),
	.S1(n336),
	.S0(n339),
	.D(\regfile[15][1] ),
	.C(\regfile[14][1] ),
	.B(\regfile[13][1] ),
	.A(\regfile[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U332 (
	.Y(n181),
	.B1(n151),
	.B0(RdData[2]),
	.A1(n361),
	.A0(N41), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U333 (
	.Y(N41),
	.S1(N13),
	.S0(N14),
	.D(n146),
	.C(n148),
	.B(n147),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U334 (
	.Y(n149),
	.S1(N12),
	.S0(n338),
	.D(REG3[2]),
	.C(REG2[2]),
	.B(REG1[2]),
	.A(REG0[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U335 (
	.Y(n147),
	.S1(N12),
	.S0(n338),
	.D(\regfile[11][2] ),
	.C(\regfile[10][2] ),
	.B(\regfile[9][2] ),
	.A(\regfile[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U336 (
	.Y(n182),
	.B1(n151),
	.B0(RdData[3]),
	.A1(n361),
	.A0(N40), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U337 (
	.Y(N40),
	.S1(N13),
	.S0(N14),
	.D(n315),
	.C(n317),
	.B(n316),
	.A(n318), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U338 (
	.Y(n318),
	.S1(N12),
	.S0(n338),
	.D(REG3[3]),
	.C(REG2[3]),
	.B(REG1[3]),
	.A(REG0[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U339 (
	.Y(n316),
	.S1(N12),
	.S0(n338),
	.D(\regfile[11][3] ),
	.C(\regfile[10][3] ),
	.B(\regfile[9][3] ),
	.A(\regfile[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U340 (
	.Y(n183),
	.B1(n151),
	.B0(RdData[4]),
	.A1(n361),
	.A0(N39), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U341 (
	.Y(N39),
	.S1(N13),
	.S0(N14),
	.D(n319),
	.C(n321),
	.B(n320),
	.A(n322), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U342 (
	.Y(n322),
	.S1(N12),
	.S0(n339),
	.D(REG3[4]),
	.C(REG2[4]),
	.B(REG1[4]),
	.A(REG0[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U343 (
	.Y(n320),
	.S1(N12),
	.S0(n338),
	.D(\regfile[11][4] ),
	.C(\regfile[10][4] ),
	.B(\regfile[9][4] ),
	.A(\regfile[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U344 (
	.Y(n184),
	.B1(n151),
	.B0(RdData[5]),
	.A1(n361),
	.A0(N38), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U345 (
	.Y(N38),
	.S1(N13),
	.S0(N14),
	.D(n323),
	.C(n325),
	.B(n324),
	.A(n326), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U346 (
	.Y(n326),
	.S1(N12),
	.S0(n339),
	.D(REG3[5]),
	.C(REG2[5]),
	.B(REG1[5]),
	.A(REG0[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U347 (
	.Y(n324),
	.S1(N12),
	.S0(n339),
	.D(\regfile[11][5] ),
	.C(\regfile[10][5] ),
	.B(\regfile[9][5] ),
	.A(\regfile[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U348 (
	.Y(n185),
	.B1(n151),
	.B0(RdData[6]),
	.A1(n361),
	.A0(N37), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U349 (
	.Y(N37),
	.S1(N13),
	.S0(N14),
	.D(n327),
	.C(n329),
	.B(n328),
	.A(n330), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U350 (
	.Y(n330),
	.S1(N12),
	.S0(n339),
	.D(REG3[6]),
	.C(REG2[6]),
	.B(REG1[6]),
	.A(REG0[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U351 (
	.Y(n328),
	.S1(N12),
	.S0(n339),
	.D(\regfile[11][6] ),
	.C(\regfile[10][6] ),
	.B(\regfile[9][6] ),
	.A(\regfile[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U352 (
	.Y(n186),
	.B1(n151),
	.B0(RdData[7]),
	.A1(n361),
	.A0(N36), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U353 (
	.Y(N36),
	.S1(N13),
	.S0(N14),
	.D(n331),
	.C(n333),
	.B(n332),
	.A(n334), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U354 (
	.Y(n334),
	.S1(N12),
	.S0(n339),
	.D(REG3[7]),
	.C(REG2[7]),
	.B(REG1[7]),
	.A(REG0[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U355 (
	.Y(n332),
	.S1(N12),
	.S0(n339),
	.D(\regfile[11][7] ),
	.C(\regfile[10][7] ),
	.B(\regfile[9][7] ),
	.A(\regfile[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U356 (
	.Y(n145),
	.S1(n336),
	.S0(n338),
	.D(REG3[1]),
	.C(REG2[1]),
	.B(REG1[1]),
	.A(REG0[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U357 (
	.Y(n140),
	.S1(n336),
	.S0(N11),
	.D(\regfile[7][0] ),
	.C(\regfile[6][0] ),
	.B(\regfile[5][0] ),
	.A(\regfile[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U358 (
	.Y(n144),
	.S1(n336),
	.S0(n338),
	.D(\regfile[7][1] ),
	.C(\regfile[6][1] ),
	.B(\regfile[5][1] ),
	.A(\regfile[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U359 (
	.Y(n148),
	.S1(N12),
	.S0(n338),
	.D(\regfile[7][2] ),
	.C(\regfile[6][2] ),
	.B(\regfile[5][2] ),
	.A(\regfile[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U360 (
	.Y(n317),
	.S1(n336),
	.S0(n338),
	.D(\regfile[7][3] ),
	.C(\regfile[6][3] ),
	.B(\regfile[5][3] ),
	.A(\regfile[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U361 (
	.Y(n321),
	.S1(N12),
	.S0(n338),
	.D(\regfile[7][4] ),
	.C(\regfile[6][4] ),
	.B(\regfile[5][4] ),
	.A(\regfile[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U362 (
	.Y(n325),
	.S1(N12),
	.S0(n339),
	.D(\regfile[7][5] ),
	.C(\regfile[6][5] ),
	.B(\regfile[5][5] ),
	.A(\regfile[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U363 (
	.Y(n329),
	.S1(N12),
	.S0(n339),
	.D(\regfile[7][6] ),
	.C(\regfile[6][6] ),
	.B(\regfile[5][6] ),
	.A(\regfile[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U364 (
	.Y(n333),
	.S1(N12),
	.S0(n339),
	.D(\regfile[7][7] ),
	.C(\regfile[6][7] ),
	.B(\regfile[5][7] ),
	.A(\regfile[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U365 (
	.Y(n138),
	.S1(n336),
	.S0(n338),
	.D(\regfile[15][0] ),
	.C(\regfile[14][0] ),
	.B(\regfile[13][0] ),
	.A(\regfile[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U366 (
	.Y(n146),
	.S1(n336),
	.S0(n338),
	.D(\regfile[15][2] ),
	.C(\regfile[14][2] ),
	.B(\regfile[13][2] ),
	.A(\regfile[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U367 (
	.Y(n315),
	.S1(n336),
	.S0(n338),
	.D(\regfile[15][3] ),
	.C(\regfile[14][3] ),
	.B(\regfile[13][3] ),
	.A(\regfile[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U368 (
	.Y(n319),
	.S1(n336),
	.S0(n338),
	.D(\regfile[15][4] ),
	.C(\regfile[14][4] ),
	.B(\regfile[13][4] ),
	.A(\regfile[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U369 (
	.Y(n323),
	.S1(n336),
	.S0(n339),
	.D(\regfile[15][5] ),
	.C(\regfile[14][5] ),
	.B(\regfile[13][5] ),
	.A(\regfile[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U370 (
	.Y(n327),
	.S1(N12),
	.S0(n339),
	.D(\regfile[15][6] ),
	.C(\regfile[14][6] ),
	.B(\regfile[13][6] ),
	.A(\regfile[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U371 (
	.Y(n331),
	.S1(N12),
	.S0(n339),
	.D(\regfile[15][7] ),
	.C(\regfile[14][7] ),
	.B(\regfile[13][7] ),
	.A(\regfile[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U372 (
	.Y(n341),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U373 (
	.Y(n178),
	.B0(n361),
	.A1(n150),
	.A0(RdData_valid), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U374 (
	.Y(n340),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U375 (
	.Y(n161),
	.B(n341),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U376 (
	.Y(n164),
	.B(n336),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U377 (
	.Y(n371),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U378 (
	.Y(n372),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U379 (
	.Y(n373),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U380 (
	.Y(n374),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module MUX_prescale (
	sel, 
	in0, 
	in1, 
	in2, 
	in3, 
	out, 
	VDD, 
	VSS);
   input [5:0] sel;
   input [7:0] in0;
   input [7:0] in1;
   input [7:0] in2;
   input [7:0] in3;
   output [7:0] out;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire FE_OFN8_n5;
   wire FE_OFN7_n6;
   wire FE_OFN6_n4;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n17;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC8_n5 (
	.Y(FE_OFN8_n5),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC7_n6 (
	.Y(FE_OFN7_n6),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX2M FE_OFC6_n4 (
	.Y(FE_OFN6_n4),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(n17),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U2 (
	.Y(n3),
	.B0(n14),
	.A2(FE_OFN7_n6),
	.A1(FE_OFN6_n4),
	.A0(FE_OFN8_n5), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U3 (
	.Y(out[1]),
	.B1(n17),
	.B0(n12),
	.A1N(n3),
	.A0N(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U4 (
	.Y(n12),
	.C1(FE_OFN7_n6),
	.C0(LTIE_LTIELO_NET),
	.B1(FE_OFN8_n5),
	.B0(LTIE_LTIELO_NET),
	.A1(FE_OFN6_n4),
	.A0(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U5 (
	.Y(out[2]),
	.B1(n17),
	.B0(n11),
	.A1N(n3),
	.A0N(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U6 (
	.Y(n11),
	.C1(FE_OFN7_n6),
	.C0(HTIE_LTIEHI_NET),
	.B1(FE_OFN8_n5),
	.B0(LTIE_LTIELO_NET),
	.A1(FE_OFN6_n4),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U7 (
	.Y(out[3]),
	.B1(n17),
	.B0(n10),
	.A1N(n3),
	.A0N(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U8 (
	.Y(n10),
	.C1(FE_OFN7_n6),
	.C0(LTIE_LTIELO_NET),
	.B1(FE_OFN8_n5),
	.B0(HTIE_LTIEHI_NET),
	.A1(FE_OFN6_n4),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U10 (
	.Y(n4),
	.D(sel[5]),
	.C(sel[3]),
	.B(sel[2]),
	.AN(sel[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U12 (
	.Y(n6),
	.D(sel[5]),
	.C(sel[4]),
	.B(sel[2]),
	.AN(sel[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U14 (
	.Y(n5),
	.D(sel[5]),
	.C(sel[4]),
	.B(sel[3]),
	.AN(sel[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n14),
	.B(sel[0]),
	.A(sel[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U16 (
	.Y(out[0]),
	.B1(n17),
	.B0(n13),
	.A1N(n3),
	.A0N(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U17 (
	.Y(n13),
	.C1(FE_OFN7_n6),
	.C0(LTIE_LTIELO_NET),
	.B1(FE_OFN8_n5),
	.B0(LTIE_LTIELO_NET),
	.A1(FE_OFN6_n4),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U18 (
	.Y(out[5]),
	.B1(n17),
	.B0(n8),
	.A1N(n3),
	.A0N(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U19 (
	.Y(n8),
	.C1(FE_OFN7_n6),
	.C0(LTIE_LTIELO_NET),
	.B1(FE_OFN8_n5),
	.B0(LTIE_LTIELO_NET),
	.A1(FE_OFN6_n4),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U20 (
	.Y(out[6]),
	.B1(n17),
	.B0(n7),
	.A1N(n3),
	.A0N(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U21 (
	.Y(n7),
	.C1(FE_OFN7_n6),
	.C0(LTIE_LTIELO_NET),
	.B1(FE_OFN8_n5),
	.B0(LTIE_LTIELO_NET),
	.A1(FE_OFN6_n4),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U22 (
	.Y(out[4]),
	.B1(n17),
	.B0(n9),
	.A1N(n3),
	.A0N(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U23 (
	.Y(n9),
	.C1(FE_OFN7_n6),
	.C0(LTIE_LTIELO_NET),
	.B1(FE_OFN8_n5),
	.B0(LTIE_LTIELO_NET),
	.A1(FE_OFN6_n4),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U24 (
	.Y(out[7]),
	.B1(n17),
	.B0(n2),
	.A1N(n3),
	.A0N(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U25 (
	.Y(n2),
	.C1(FE_OFN7_n6),
	.C0(LTIE_LTIELO_NET),
	.B1(FE_OFN8_n5),
	.B0(LTIE_LTIELO_NET),
	.A1(FE_OFN6_n4),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clock_divider_test_0 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	CLK_UART_M__L10_N0, 
	CLK_UART_M__L5_N0, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input CLK_UART_M__L10_N0;
   input CLK_UART_M__L5_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN9_o_div_clk_reg__Exclude_0_NET;
   wire o_div_clk_reg__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire o_div_clk_reg;
   wire flag;
   wire N9;
   wire N12;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire [7:0] half_toggle;
   wire [7:0] half_toggle_p1;
   wire [6:0] counter;

//   assign test_so = n55 ;

   // Module instantiations
   DLY3X1M FE_PHC9_o_div_clk_reg__Exclude_0_NET (
	.Y(FE_PHN9_o_div_clk_reg__Exclude_0_NET),
	.A(o_div_clk_reg__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M o_div_clk_reg__Exclude_0 (
	.Y(o_div_clk_reg__Exclude_0_NET),
	.A(o_div_clk_reg), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M flag_reg (
	.SI(counter[6]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(flag),
	.D(n34),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M o_div_clk_reg_reg (
	.SI(flag),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(o_div_clk_reg),
	.D(n33),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(n37),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[6]),
	.D(N42),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[5]),
	.D(N41),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(n36),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[4]),
	.D(N40),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[0]),
	.D(N36),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(counter[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[1]),
	.D(N37),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[3]),
	.D(N39),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[2]),
	.D(N38),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n52),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U6 (
	.Y(n34),
	.B(n26),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(n28),
	.B(n54),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(N37),
	.B(n52),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(N38),
	.B(n52),
	.A(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U17 (
	.Y(N39),
	.B(n52),
	.A(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U18 (
	.Y(N40),
	.B(n52),
	.A(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U19 (
	.Y(N41),
	.B(n52),
	.A(N21), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n53),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n51),
	.A(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n45),
	.A(half_toggle_p1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n46),
	.A(half_toggle_p1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n47),
	.A(half_toggle_p1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n48),
	.A(half_toggle_p1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n22),
	.A(half_toggle[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n23),
	.A(half_toggle[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n24),
	.A(half_toggle[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n25),
	.A(half_toggle[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U30 (
	.Y(n27),
	.C0(n53),
	.B0(n29),
	.A1N(N9),
	.A0(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U31 (
	.Y(n33),
	.B1(test_so),
	.B0(n27),
	.A2(n52),
	.A1(o_div_clk_reg__Exclude_0_NET),
	.A0(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(test_so),
	.A(FE_PHN9_o_div_clk_reg__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(half_toggle[0]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U34 (
	.Y(n29),
	.B(i_div_ratio[0]),
	.AN(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U35 (
	.Y(n30),
	.B1(N9),
	.B0(flag),
	.A1(n54),
	.A0(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U36 (
	.Y(N42),
	.B(n52),
	.A(N22), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U37 (
	.Y(N36),
	.B(n52),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n49),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n35),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n36),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U41 (
	.Y(n26),
	.B0(HTIE_LTIEHI_NET),
	.A1N(n32),
	.A0N(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U42 (
	.Y(n31),
	.C(i_div_ratio[2]),
	.B(i_div_ratio[3]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U43 (
	.Y(n32),
	.D(i_div_ratio[4]),
	.C(i_div_ratio[5]),
	.B(i_div_ratio[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n50),
	.A(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n37),
	.A(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n54),
	.A(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U47 (
	.Y(o_div_clk),
	.S0(n53),
	.B(o_div_clk_reg),
	.A(CLK_UART_M__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U48 (
	.Y(n1),
	.B(half_toggle[0]),
	.AN(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U49 (
	.Y(half_toggle[1]),
	.B0(n1),
	.A1N(i_div_ratio[2]),
	.A0N(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U50 (
	.Y(n2),
	.B(i_div_ratio[3]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U51 (
	.Y(half_toggle[2]),
	.B0(n2),
	.A1N(i_div_ratio[3]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U52 (
	.Y(n3),
	.B(i_div_ratio[4]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U53 (
	.Y(half_toggle[3]),
	.B0(n3),
	.A1N(i_div_ratio[4]),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U54 (
	.Y(n4),
	.B(i_div_ratio[5]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U55 (
	.Y(half_toggle[4]),
	.B0(n4),
	.A1N(i_div_ratio[5]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U56 (
	.Y(half_toggle[5]),
	.B(n4),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U57 (
	.Y(half_toggle[7]),
	.C(n4),
	.B(i_div_ratio[7]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U58 (
	.Y(n5),
	.B0(i_div_ratio[7]),
	.A1(n4),
	.A0(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U59 (
	.Y(half_toggle[6]),
	.B(n5),
	.AN(half_toggle[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U60 (
	.Y(n6),
	.B0(counter[0]),
	.A1N(n49),
	.A0N(half_toggle[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U61 (
	.Y(n7),
	.C1(n49),
	.C0(half_toggle[1]),
	.B1(half_toggle[0]),
	.B0(n6),
	.A1(n35),
	.A0(half_toggle[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U62 (
	.Y(n8),
	.C0(n7),
	.B1(n22),
	.B0(counter[2]),
	.A1(n23),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U63 (
	.Y(n9),
	.C0(n8),
	.B1(n36),
	.B0(half_toggle[3]),
	.A1(n50),
	.A0(half_toggle[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U64 (
	.Y(n10),
	.C0(n9),
	.B1(n24),
	.B0(counter[4]),
	.A1(n25),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U65 (
	.Y(n11),
	.C0(n10),
	.B1(n37),
	.B0(half_toggle[5]),
	.A1(n51),
	.A0(half_toggle[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U66 (
	.Y(n12),
	.B0(n11),
	.A1N(n51),
	.A0N(half_toggle[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(N9),
	.B(n12),
	.A(half_toggle[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U68 (
	.Y(n38),
	.B0(counter[0]),
	.A1N(n49),
	.A0N(half_toggle_p1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U69 (
	.Y(n39),
	.C1(n49),
	.C0(half_toggle_p1[1]),
	.B1(half_toggle_p1[0]),
	.B0(n38),
	.A1(n35),
	.A0(half_toggle_p1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U70 (
	.Y(n40),
	.C0(n39),
	.B1(n45),
	.B0(counter[2]),
	.A1(n46),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U71 (
	.Y(n41),
	.C0(n40),
	.B1(n36),
	.B0(half_toggle_p1[3]),
	.A1(n50),
	.A0(half_toggle_p1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U72 (
	.Y(n42),
	.C0(n41),
	.B1(n47),
	.B0(counter[4]),
	.A1(n48),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U73 (
	.Y(n43),
	.C0(n42),
	.B1(n37),
	.B0(half_toggle_p1[5]),
	.A1(n51),
	.A0(half_toggle_p1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U74 (
	.Y(n44),
	.B0(n43),
	.A1N(n51),
	.A0N(half_toggle_p1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(N12),
	.B(n44),
	.A(half_toggle_p1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   clock_divider_0_DW01_inc_0 add_39 (
	.A({ counter[6],
		counter[5],
		counter[4],
		counter[3],
		counter[2],
		counter[1],
		counter[0] }),
	.SUM({ N22,
		N21,
		N20,
		N19,
		N18,
		N17,
		N16 }), 
	.VDD(VDD), 
	.VSS(VSS));
   clock_divider_0_DW01_inc_1 add_18 (
	.A({ half_toggle[7],
		half_toggle[6],
		half_toggle[5],
		half_toggle[4],
		half_toggle[3],
		half_toggle[2],
		half_toggle[1],
		half_toggle[0] }),
	.SUM({ half_toggle_p1[7],
		half_toggle_p1[6],
		half_toggle_p1[5],
		half_toggle_p1[4],
		half_toggle_p1[3],
		half_toggle_p1[2],
		half_toggle_p1[1],
		half_toggle_p1[0] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clock_divider_0_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [6:0] A;
   output [6:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [6:2] carry;

   // Module instantiations
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[6]),
	.B(A[6]),
	.A(carry[6]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clock_divider_0_DW01_inc_1 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clock_divider_test_1 (
	i_ref_clk, 
	i_rst_n, 
	i_clk_en, 
	i_div_ratio, 
	o_div_clk, 
	test_si, 
	test_so, 
	test_se, 
	CLK_UART_M__L10_N0, 
	CLK_UART_M__L5_N0, 
	VDD, 
	VSS);
   input i_ref_clk;
   input i_rst_n;
   input i_clk_en;
   input [7:0] i_div_ratio;
   output o_div_clk;
   input test_si;
   output test_so;
   input test_se;
   input CLK_UART_M__L10_N0;
   input CLK_UART_M__L5_N0;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_PHN8_o_div_clk_reg__Exclude_0_NET;
   wire o_div_clk_reg__Exclude_0_NET;
   wire HTIE_LTIEHI_NET;
   wire o_div_clk_reg;
   wire flag;
   wire N9;
   wire N12;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N21;
   wire N22;
   wire N36;
   wire N37;
   wire N38;
   wire N39;
   wire N40;
   wire N41;
   wire N42;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire [7:0] half_toggle;
   wire [7:0] half_toggle_p1;
   wire [6:0] counter;

//   assign test_so = n54 ;

   // Module instantiations
   DLY3X1M FE_PHC8_o_div_clk_reg__Exclude_0_NET (
	.Y(FE_PHN8_o_div_clk_reg__Exclude_0_NET),
	.A(o_div_clk_reg__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   BUFX8M o_div_clk_reg__Exclude_0 (
	.Y(o_div_clk_reg__Exclude_0_NET),
	.A(o_div_clk_reg), 
	.VDD(VDD), 
	.VSS(VSS));
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M flag_reg (
	.SI(counter[6]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(flag),
	.D(n56),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M o_div_clk_reg_reg (
	.SI(flag),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(o_div_clk_reg),
	.D(n57),
	.CK(i_ref_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[6]  (
	.SI(n37),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[6]),
	.D(N42),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[5]  (
	.SI(counter[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[5]),
	.D(N41),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[4]  (
	.SI(n36),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[4]),
	.D(N40),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[0]),
	.D(N36),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(counter[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[1]),
	.D(N37),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(counter[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[3]),
	.D(N39),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(counter[2]),
	.D(N38),
	.CK(CLK_UART_M__L10_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n52),
	.A(n63), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X2M U6 (
	.Y(n63),
	.C0(n55),
	.B0(n61),
	.A1N(N9),
	.A0(i_div_ratio[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(half_toggle[0]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(N37),
	.B(n52),
	.A(N17), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(N38),
	.B(n52),
	.A(N18), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U17 (
	.Y(N39),
	.B(n52),
	.A(N19), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U18 (
	.Y(N40),
	.B(n52),
	.A(N20), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U19 (
	.Y(N41),
	.B(n52),
	.A(N21), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U20 (
	.Y(n56),
	.B(n64),
	.A(n62), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U21 (
	.Y(n62),
	.B(n53),
	.A(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n55),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n51),
	.A(counter[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n45),
	.A(half_toggle_p1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U25 (
	.Y(n46),
	.A(half_toggle_p1[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n47),
	.A(half_toggle_p1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n48),
	.A(half_toggle_p1[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n25),
	.A(half_toggle[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n24),
	.A(half_toggle[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U30 (
	.Y(n23),
	.A(half_toggle[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(n22),
	.A(half_toggle[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U32 (
	.Y(n57),
	.B1(test_so),
	.B0(n63),
	.A2(n52),
	.A1(o_div_clk_reg__Exclude_0_NET),
	.A0(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(test_so),
	.A(FE_PHN8_o_div_clk_reg__Exclude_0_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U34 (
	.Y(n61),
	.B(i_div_ratio[0]),
	.AN(n60), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U35 (
	.Y(n60),
	.B1(N9),
	.B0(flag),
	.A1(n53),
	.A0(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U36 (
	.Y(N42),
	.B(n52),
	.A(N22), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U37 (
	.Y(N36),
	.B(n52),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U38 (
	.Y(n49),
	.A(counter[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n35),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n36),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U41 (
	.Y(n64),
	.B0(HTIE_LTIEHI_NET),
	.A1N(n58),
	.A0N(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U42 (
	.Y(n58),
	.D(i_div_ratio[4]),
	.C(i_div_ratio[5]),
	.B(i_div_ratio[6]),
	.A(i_div_ratio[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U43 (
	.Y(n59),
	.C(i_div_ratio[2]),
	.B(i_div_ratio[3]),
	.A(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n50),
	.A(counter[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U45 (
	.Y(n37),
	.A(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n53),
	.A(flag), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U47 (
	.Y(o_div_clk),
	.S0(n55),
	.B(o_div_clk_reg),
	.A(CLK_UART_M__L5_N0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U48 (
	.Y(n1),
	.B(half_toggle[0]),
	.AN(i_div_ratio[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U49 (
	.Y(half_toggle[1]),
	.B0(n1),
	.A1N(i_div_ratio[2]),
	.A0N(i_div_ratio[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U50 (
	.Y(n2),
	.B(i_div_ratio[3]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U51 (
	.Y(half_toggle[2]),
	.B0(n2),
	.A1N(i_div_ratio[3]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U52 (
	.Y(n3),
	.B(i_div_ratio[4]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U53 (
	.Y(half_toggle[3]),
	.B0(n3),
	.A1N(i_div_ratio[4]),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U54 (
	.Y(n4),
	.B(i_div_ratio[5]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U55 (
	.Y(half_toggle[4]),
	.B0(n4),
	.A1N(i_div_ratio[5]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U56 (
	.Y(half_toggle[5]),
	.B(n4),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U57 (
	.Y(half_toggle[7]),
	.C(n4),
	.B(i_div_ratio[7]),
	.A(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U58 (
	.Y(n5),
	.B0(i_div_ratio[7]),
	.A1(n4),
	.A0(i_div_ratio[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U59 (
	.Y(half_toggle[6]),
	.B(n5),
	.AN(half_toggle[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U60 (
	.Y(n6),
	.B0(counter[0]),
	.A1N(n49),
	.A0N(half_toggle[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U61 (
	.Y(n7),
	.C1(n49),
	.C0(half_toggle[1]),
	.B1(half_toggle[0]),
	.B0(n6),
	.A1(n35),
	.A0(half_toggle[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U62 (
	.Y(n8),
	.C0(n7),
	.B1(n25),
	.B0(counter[2]),
	.A1(n24),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U63 (
	.Y(n9),
	.C0(n8),
	.B1(n36),
	.B0(half_toggle[3]),
	.A1(n50),
	.A0(half_toggle[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U64 (
	.Y(n10),
	.C0(n9),
	.B1(n23),
	.B0(counter[4]),
	.A1(n22),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U65 (
	.Y(n11),
	.C0(n10),
	.B1(n37),
	.B0(half_toggle[5]),
	.A1(n51),
	.A0(half_toggle[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U66 (
	.Y(n12),
	.B0(n11),
	.A1N(n51),
	.A0N(half_toggle[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(N9),
	.B(n12),
	.A(half_toggle[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U68 (
	.Y(n38),
	.B0(counter[0]),
	.A1N(n49),
	.A0N(half_toggle_p1[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U69 (
	.Y(n39),
	.C1(n49),
	.C0(half_toggle_p1[1]),
	.B1(half_toggle_p1[0]),
	.B0(n38),
	.A1(n35),
	.A0(half_toggle_p1[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U70 (
	.Y(n40),
	.C0(n39),
	.B1(n45),
	.B0(counter[2]),
	.A1(n46),
	.A0(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U71 (
	.Y(n41),
	.C0(n40),
	.B1(n36),
	.B0(half_toggle_p1[3]),
	.A1(n50),
	.A0(half_toggle_p1[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U72 (
	.Y(n42),
	.C0(n41),
	.B1(n47),
	.B0(counter[4]),
	.A1(n48),
	.A0(counter[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U73 (
	.Y(n43),
	.C0(n42),
	.B1(n37),
	.B0(half_toggle_p1[5]),
	.A1(n51),
	.A0(half_toggle_p1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U74 (
	.Y(n44),
	.B0(n43),
	.A1N(n51),
	.A0N(half_toggle_p1[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(N12),
	.B(n44),
	.A(half_toggle_p1[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   clock_divider_1_DW01_inc_0 add_39 (
	.A({ counter[6],
		counter[5],
		counter[4],
		counter[3],
		counter[2],
		counter[1],
		counter[0] }),
	.SUM({ N22,
		N21,
		N20,
		N19,
		N18,
		N17,
		N16 }), 
	.VDD(VDD), 
	.VSS(VSS));
   clock_divider_1_DW01_inc_1 add_18 (
	.A({ half_toggle[7],
		half_toggle[6],
		half_toggle[5],
		half_toggle[4],
		half_toggle[3],
		half_toggle[2],
		half_toggle[1],
		half_toggle[0] }),
	.SUM({ half_toggle_p1[7],
		half_toggle_p1[6],
		half_toggle_p1[5],
		half_toggle_p1[4],
		half_toggle_p1[3],
		half_toggle_p1[2],
		half_toggle_p1[1],
		half_toggle_p1[0] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clock_divider_1_DW01_inc_0 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [6:0] A;
   output [6:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [6:2] carry;

   // Module instantiations
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[6]),
	.B(A[6]),
	.A(carry[6]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module clock_divider_1_DW01_inc_1 (
	A, 
	SUM, 
	VDD, 
	VSS);
   input [7:0] A;
   output [7:0] SUM;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [7:2] carry;

   // Module instantiations
   ADDHX1M U1_1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.B(A[0]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.B(carry[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.B(carry[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.B(carry[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.B(carry[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U1_1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.B(carry[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U1 (
	.Y(SUM[0]),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[7]),
	.B(A[7]),
	.A(carry[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module PULSE_GEN_test_1 (
	CLK, 
	RST_n, 
	LVL_SIG, 
	pulse_out, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK;
   input RST_n;
   input LVL_SIG;
   output pulse_out;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire LVL_SIG_reg;

   assign test_so = LVL_SIG_reg ;

   // Module instantiations
   SDFFRQX2M LVL_SIG_reg_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_n),
	.Q(LVL_SIG_reg),
	.D(LVL_SIG),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U4 (
	.Y(pulse_out),
	.B(LVL_SIG_reg),
	.AN(LVL_SIG), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_test_1 (
	CLK, 
	RST, 
	A, 
	B, 
	ALU_FUN, 
	Enable, 
	valid_data, 
	ALU_OUT, 
	test_si, 
	test_se, 
	FE_OFN0_RST_SYNC_1_mux, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] A;
   input [7:0] B;
   input [3:0] ALU_FUN;
   input Enable;
   output valid_data;
   output [15:0] ALU_OUT;
   input test_si;
   input test_se;
   input FE_OFN0_RST_SYNC_1_mux;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN5_n50;
   wire N92;
   wire N93;
   wire N94;
   wire N95;
   wire N96;
   wire N97;
   wire N98;
   wire N99;
   wire N100;
   wire N101;
   wire N102;
   wire N103;
   wire N104;
   wire N105;
   wire N106;
   wire N107;
   wire N108;
   wire N109;
   wire N110;
   wire N111;
   wire N112;
   wire N113;
   wire N114;
   wire N115;
   wire N116;
   wire N117;
   wire N118;
   wire N119;
   wire N120;
   wire N121;
   wire N122;
   wire N123;
   wire N124;
   wire N125;
   wire N126;
   wire N127;
   wire N128;
   wire N129;
   wire N130;
   wire N131;
   wire N132;
   wire N133;
   wire N166;
   wire N167;
   wire N168;
   wire N185;
   wire N186;
   wire N187;
   wire N188;
   wire N189;
   wire N190;
   wire N191;
   wire N192;
   wire N193;
   wire N194;
   wire N195;
   wire N196;
   wire N197;
   wire N198;
   wire N199;
   wire N200;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n82;
   wire n83;
   wire n84;
   wire n85;
   wire n86;
   wire n87;
   wire n88;
   wire n89;
   wire n90;
   wire n91;
   wire n92;
   wire n93;
   wire n94;
   wire n95;
   wire n96;
   wire n97;
   wire n98;
   wire n99;
   wire n100;
   wire n101;
   wire n102;
   wire n103;
   wire n104;
   wire n105;
   wire n106;
   wire n107;
   wire n108;
   wire n109;
   wire n110;
   wire n111;
   wire n112;
   wire n113;
   wire n114;
   wire n115;
   wire n116;
   wire n117;
   wire n118;
   wire n119;
   wire n120;
   wire n121;
   wire n122;
   wire n123;
   wire n124;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n125;
   wire n126;
   wire n127;
   wire n128;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;

   // Module instantiations
   BUFX2M FE_OFC5_n50 (
	.Y(FE_OFN5_n50),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[7]  (
	.SI(ALU_OUT[6]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[7]),
	.D(N192),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[6]  (
	.SI(ALU_OUT[5]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[6]),
	.D(N191),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[5]  (
	.SI(ALU_OUT[4]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[5]),
	.D(N190),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[4]  (
	.SI(ALU_OUT[3]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[4]),
	.D(N189),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[3]  (
	.SI(ALU_OUT[2]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[3]),
	.D(N188),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \ALU_OUT_reg[2]  (
	.SI(ALU_OUT[1]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[2]),
	.D(N187),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \ALU_OUT_reg[1]  (
	.SI(ALU_OUT[0]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[1]),
	.D(N186),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRHQX1M \ALU_OUT_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[0]),
	.D(N185),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[15]  (
	.SI(ALU_OUT[14]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[15]),
	.D(N200),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[14]  (
	.SI(ALU_OUT[13]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[14]),
	.D(N199),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[13]  (
	.SI(ALU_OUT[12]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[13]),
	.D(N198),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[12]  (
	.SI(ALU_OUT[11]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[12]),
	.D(N197),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[11]  (
	.SI(ALU_OUT[10]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[11]),
	.D(N196),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[10]  (
	.SI(ALU_OUT[9]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[10]),
	.D(N195),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[9]  (
	.SI(ALU_OUT[8]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(ALU_OUT[9]),
	.D(N194),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \ALU_OUT_reg[8]  (
	.SI(ALU_OUT[7]),
	.SE(test_se),
	.RN(RST),
	.Q(ALU_OUT[8]),
	.D(N193),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX1M valid_data_reg (
	.SI(ALU_OUT[15]),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(valid_data),
	.D(Enable),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U24 (
	.Y(n58),
	.B0(n118),
	.A1N(n122),
	.A0N(n147), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U25 (
	.Y(n67),
	.B0(n118),
	.A1N(n116),
	.A0N(n117), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U26 (
	.Y(n54),
	.B(n144),
	.AN(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U27 (
	.Y(n143),
	.A(ALU_FUN[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U28 (
	.Y(n62),
	.B(n122),
	.A(n116), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n56),
	.B(n122),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U31 (
	.Y(n57),
	.B(n144),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n144),
	.A(n117), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U33 (
	.Y(n145),
	.A(n109), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(n147),
	.A(n124), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U35 (
	.Y(n48),
	.B(n142),
	.AN(FE_OFN5_n50), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U36 (
	.Y(N194),
	.B0(n49),
	.A1N(n48),
	.A0N(N119), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U37 (
	.Y(N195),
	.B0(n49),
	.A1N(n48),
	.A0N(N120), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U38 (
	.Y(N196),
	.B0(n49),
	.A1N(n48),
	.A0N(N121), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U39 (
	.Y(N197),
	.B0(n49),
	.A1N(n48),
	.A0N(N122), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U40 (
	.Y(N198),
	.B0(n49),
	.A1N(n48),
	.A0N(N123), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U41 (
	.Y(N199),
	.B0(n49),
	.A1N(n48),
	.A0N(N124), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U42 (
	.Y(N200),
	.B0(n49),
	.A1N(n48),
	.A0N(N125), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3BX4M U43 (
	.Y(n68),
	.C(ALU_FUN[2]),
	.B(n146),
	.AN(n122), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U44 (
	.Y(n50),
	.C(n146),
	.B(ALU_FUN[2]),
	.A(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U45 (
	.Y(n123),
	.B(ALU_FUN[1]),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U46 (
	.Y(n66),
	.C(ALU_FUN[3]),
	.B(n143),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U47 (
	.Y(n53),
	.C(ALU_FUN[3]),
	.B(n143),
	.A(n147), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U48 (
	.Y(n124),
	.B(ALU_FUN[1]),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U49 (
	.Y(n122),
	.B(ALU_FUN[3]),
	.A(n143), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U50 (
	.Y(n117),
	.B(ALU_FUN[0]),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U51 (
	.Y(n109),
	.C(n116),
	.B(ALU_FUN[0]),
	.A(ALU_FUN[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U52 (
	.Y(n146),
	.A(ALU_FUN[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U53 (
	.Y(n118),
	.C(ALU_FUN[3]),
	.B(ALU_FUN[0]),
	.A(n123), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U54 (
	.Y(n116),
	.B(n146),
	.A(ALU_FUN[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U55 (
	.Y(n108),
	.D(n143),
	.C(ALU_FUN[3]),
	.B(n116),
	.A(N168), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U56 (
	.Y(n49),
	.B(n141),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U57 (
	.Y(N187),
	.B0(n142),
	.A2(n95),
	.A1(n94),
	.A0(n93), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U58 (
	.Y(n93),
	.B1(n54),
	.B0(N94),
	.A1(n56),
	.A0(N103), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U59 (
	.Y(n95),
	.C0(n96),
	.B1(n156),
	.B0(n57),
	.A1(n145),
	.A0(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U60 (
	.Y(n94),
	.C1(n68),
	.C0(N128),
	.B1(n62),
	.B0(A[2]),
	.A1(FE_OFN5_n50),
	.A0(N112), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U61 (
	.Y(N188),
	.B0(n142),
	.A2(n89),
	.A1(n88),
	.A0(n87), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U62 (
	.Y(n87),
	.B1(n54),
	.B0(N95),
	.A1(n56),
	.A0(N104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U63 (
	.Y(n89),
	.C0(n90),
	.B1(n155),
	.B0(n57),
	.A1(n145),
	.A0(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U64 (
	.Y(n88),
	.C1(n68),
	.C0(N129),
	.B1(n62),
	.B0(A[3]),
	.A1(FE_OFN5_n50),
	.A0(N113), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U65 (
	.Y(N189),
	.B0(n142),
	.A2(n83),
	.A1(n82),
	.A0(n81), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U66 (
	.Y(n81),
	.B1(n54),
	.B0(N96),
	.A1(n56),
	.A0(N105), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U67 (
	.Y(n83),
	.C0(n84),
	.B1(n154),
	.B0(n57),
	.A1(A[5]),
	.A0(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U68 (
	.Y(n82),
	.C1(n68),
	.C0(N130),
	.B1(n62),
	.B0(A[4]),
	.A1(FE_OFN5_n50),
	.A0(N114), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U69 (
	.Y(N190),
	.B0(n142),
	.A2(n77),
	.A1(n76),
	.A0(n75), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U70 (
	.Y(n75),
	.B1(n54),
	.B0(N97),
	.A1(n56),
	.A0(N106), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U71 (
	.Y(n77),
	.C0(n78),
	.B1(n153),
	.B0(n57),
	.A1(A[6]),
	.A0(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U72 (
	.Y(n76),
	.C1(n68),
	.C0(N131),
	.B1(n62),
	.B0(A[5]),
	.A1(FE_OFN5_n50),
	.A0(N115), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U73 (
	.Y(N191),
	.B0(n142),
	.A2(n71),
	.A1(n70),
	.A0(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U74 (
	.Y(n69),
	.B1(n54),
	.B0(N98),
	.A1(n56),
	.A0(N107), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U75 (
	.Y(n71),
	.C0(n72),
	.B1(n152),
	.B0(n57),
	.A1(A[7]),
	.A0(n145), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U76 (
	.Y(n70),
	.C1(n68),
	.C0(N132),
	.B1(A[6]),
	.B0(n62),
	.A1(FE_OFN5_n50),
	.A0(N116), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U77 (
	.Y(N192),
	.B0(n142),
	.A2(n61),
	.A1(n60),
	.A0(n59), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U78 (
	.Y(n60),
	.B1(FE_OFN5_n50),
	.B0(N117),
	.A1(n68),
	.A0(N133), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U79 (
	.Y(n59),
	.B1(n54),
	.B0(N99),
	.A1(n56),
	.A0(N108), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U80 (
	.Y(n61),
	.C0(n63),
	.B1(A[7]),
	.B0(n62),
	.A1(n151),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U81 (
	.Y(N185),
	.B0(n142),
	.A2(n112),
	.A1(n111),
	.A0(n110), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U82 (
	.Y(n110),
	.B1(n54),
	.B0(N92),
	.A1(n56),
	.A0(N101), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U83 (
	.Y(n112),
	.C0(n114),
	.B0(n113),
	.A1(n158),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X4M U84 (
	.Y(n111),
	.C1(n68),
	.C0(N126),
	.B1(n62),
	.B0(A[0]),
	.A1(FE_OFN5_n50),
	.A0(N110), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U85 (
	.Y(N186),
	.B0(n142),
	.A2(n101),
	.A1(n100),
	.A0(n99), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U86 (
	.Y(n101),
	.C0(n103),
	.B0(n102),
	.A1(n145),
	.A0(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U87 (
	.Y(n100),
	.C1(n62),
	.C0(A[1]),
	.B1(n157),
	.B0(n57),
	.A1(n68),
	.A0(N127), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI222X1M U88 (
	.Y(n99),
	.C1(n56),
	.C0(N102),
	.B1(FE_OFN5_n50),
	.B0(N111),
	.A1(n54),
	.A0(N93), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U89 (
	.Y(n142),
	.A(Enable), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U90 (
	.Y(N193),
	.B0(n142),
	.A1(n52),
	.A0(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U91 (
	.Y(n51),
	.B0(n141),
	.A1(n54),
	.A0(N100), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2XLM U92 (
	.Y(n52),
	.B1(FE_OFN5_n50),
	.B0(N118),
	.A1N(n53),
	.A0N(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U93 (
	.Y(n72),
	.C1(n153),
	.C0(n53),
	.B1(n74),
	.B0(B[6]),
	.A1(n140),
	.A0(n73), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U94 (
	.Y(n74),
	.C0(n57),
	.B1(n152),
	.B0(n58),
	.A1(n66),
	.A0(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U95 (
	.Y(n73),
	.C0(n62),
	.B1(n67),
	.B0(A[6]),
	.A1(n152),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U96 (
	.Y(n138),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U97 (
	.Y(n141),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U98 (
	.Y(n55),
	.C0(n58),
	.B0(n57),
	.A1(n56),
	.A0(N109), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U99 (
	.Y(N167),
	.A(n134), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U100 (
	.Y(n140),
	.A(B[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U102 (
	.Y(n157),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U103 (
	.Y(n158),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U104 (
	.Y(n152),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U105 (
	.Y(n151),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U106 (
	.Y(n155),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U107 (
	.Y(n156),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n153),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U109 (
	.Y(n154),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U110 (
	.Y(n96),
	.C1(n157),
	.C0(n53),
	.B1(n98),
	.B0(B[2]),
	.A1(n137),
	.A0(n97), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U111 (
	.Y(n98),
	.C0(n57),
	.B1(n156),
	.B0(n58),
	.A1(n66),
	.A0(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U112 (
	.Y(n97),
	.C0(n62),
	.B1(n67),
	.B0(A[2]),
	.A1(n156),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U113 (
	.Y(n90),
	.C1(n156),
	.C0(n53),
	.B1(n92),
	.B0(B[3]),
	.A1(n139),
	.A0(n91), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U114 (
	.Y(n92),
	.C0(n57),
	.B1(n155),
	.B0(n58),
	.A1(n66),
	.A0(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U115 (
	.Y(n91),
	.C0(n62),
	.B1(n67),
	.B0(A[3]),
	.A1(n155),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U116 (
	.Y(n84),
	.C1(n155),
	.C0(n53),
	.B1(n86),
	.B0(B[4]),
	.A1(n150),
	.A0(n85), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U117 (
	.Y(n150),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U118 (
	.Y(n86),
	.C0(n57),
	.B1(n154),
	.B0(n58),
	.A1(n66),
	.A0(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U119 (
	.Y(n85),
	.C0(n62),
	.B1(n67),
	.B0(A[4]),
	.A1(n154),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U120 (
	.Y(n78),
	.C1(n154),
	.C0(n53),
	.B1(n80),
	.B0(B[5]),
	.A1(n149),
	.A0(n79), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U121 (
	.Y(n149),
	.A(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U122 (
	.Y(n80),
	.C0(n57),
	.B1(n153),
	.B0(n58),
	.A1(n66),
	.A0(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U123 (
	.Y(n79),
	.C0(n62),
	.B1(n67),
	.B0(A[5]),
	.A1(n153),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI222X1M U124 (
	.Y(n63),
	.C1(n152),
	.C0(n53),
	.B1(n65),
	.B0(B[7]),
	.A1(n148),
	.A0(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U125 (
	.Y(n148),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U126 (
	.Y(n65),
	.C0(n57),
	.B1(n151),
	.B0(n58),
	.A1(A[7]),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U127 (
	.Y(n64),
	.C0(n62),
	.B1(n67),
	.B0(A[7]),
	.A1(n151),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U128 (
	.Y(n136),
	.A(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U129 (
	.Y(n114),
	.B1(n157),
	.B0(n109),
	.A1N(B[0]),
	.A0(n115), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U130 (
	.Y(n115),
	.C0(n62),
	.B1(n67),
	.B0(A[0]),
	.A1(n158),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U131 (
	.Y(n103),
	.B1(n158),
	.B0(n53),
	.A1N(B[1]),
	.A0(n104), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U132 (
	.Y(n104),
	.C0(n62),
	.B1(n67),
	.B0(A[1]),
	.A1(n157),
	.A0(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U133 (
	.Y(n113),
	.B0(n120),
	.A1(n119),
	.A0(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U134 (
	.Y(n120),
	.B0(n108),
	.A2(n121),
	.A1(ALU_FUN[3]),
	.A0(N166), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U135 (
	.Y(n119),
	.C0(n57),
	.B1(n158),
	.B0(n58),
	.A1(n66),
	.A0(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U136 (
	.Y(n121),
	.C(ALU_FUN[0]),
	.B(ALU_FUN[2]),
	.A(n146), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U137 (
	.Y(n102),
	.B0(n106),
	.A1(n105),
	.A0(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U138 (
	.Y(n106),
	.B0(n108),
	.A2(n107),
	.A1(ALU_FUN[3]),
	.A0(N167), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI221XLM U139 (
	.Y(n105),
	.C0(n57),
	.B1(n157),
	.B0(n58),
	.A1(n66),
	.A0(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U140 (
	.Y(n107),
	.C(n146),
	.B(ALU_FUN[2]),
	.A(n143), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U149 (
	.Y(n135),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U150 (
	.Y(n137),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U151 (
	.Y(n139),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U152 (
	.Y(n131),
	.B(B[7]),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U153 (
	.Y(n47),
	.B(A[4]),
	.AN(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U154 (
	.Y(n36),
	.B(B[4]),
	.AN(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U155 (
	.Y(n126),
	.B(n36),
	.A(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U156 (
	.Y(n44),
	.B(A[3]),
	.A(n139), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U157 (
	.Y(n35),
	.B(A[2]),
	.A(n137), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U158 (
	.Y(n32),
	.B(A[0]),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U159 (
	.Y(n46),
	.B(n137),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U160 (
	.Y(n41),
	.B(n46),
	.AN(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U161 (
	.Y(n33),
	.B0(B[1]),
	.A1(n157),
	.A0(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U162 (
	.Y(n34),
	.C0(n33),
	.B0(n41),
	.A1(n136),
	.A0(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U163 (
	.Y(n45),
	.B(n139),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U164 (
	.Y(n37),
	.B0(n45),
	.A2(n34),
	.A1(n35),
	.A0(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U165 (
	.Y(n129),
	.B(B[5]),
	.AN(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X1M U166 (
	.Y(n38),
	.C0(n129),
	.B0(n36),
	.A1(n37),
	.A0(n126), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U167 (
	.Y(n125),
	.B(A[5]),
	.AN(B[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U168 (
	.Y(n128),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U169 (
	.Y(n39),
	.B1(n152),
	.B0(B[6]),
	.A2(n128),
	.A1(n125),
	.A0(n38), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U170 (
	.Y(n132),
	.B(n151),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U171 (
	.Y(N168),
	.B0(n132),
	.A1(n39),
	.A0(n131), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U172 (
	.Y(n42),
	.B(n135),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U173 (
	.Y(n40),
	.B0(B[1]),
	.A1(n157),
	.A0(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X1M U174 (
	.Y(n43),
	.C0(n40),
	.B0(n41),
	.A1(n157),
	.A0(n42), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X1M U175 (
	.Y(n127),
	.B0(n44),
	.A2(n45),
	.A1(n46),
	.A0(n138), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X1M U176 (
	.Y(n130),
	.C0(n47),
	.B0(n125),
	.A1N(n127),
	.A0(n126), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U177 (
	.Y(n133),
	.B1(n140),
	.B0(A[6]),
	.A2(n128),
	.A1(n129),
	.A0(n130), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U178 (
	.Y(n134),
	.B0(n131),
	.A1N(n133),
	.A0(n132), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U179 (
	.Y(N166),
	.B(N167),
	.A(N168), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW_div_uns_0 div_29 (
	.a({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.b({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.quotient({ N133,
		N132,
		N131,
		N130,
		N129,
		N128,
		N127,
		N126 }),
	.n148(n148),
	.n158(n158),
	.n157(n157),
	.n140(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_sub_0 sub_27 (
	.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.CI(1'b0),
	.DIFF({ N109,
		N108,
		N107,
		N106,
		N105,
		N104,
		N103,
		N102,
		N101 }),
	.n135(n135),
	.n137(n137),
	.n139(n139),
	.n148(n148),
	.n150(n150),
	.n149(n149),
	.n158(n158),
	.n140(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_add_0 add_26 (
	.A({ 1'b0,
		A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ 1'b0,
		B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.CI(1'b0),
	.SUM({ N100,
		N99,
		N98,
		N97,
		N96,
		N95,
		N94,
		N93,
		N92 }), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW02_mult_0 mult_28 (
	.A({ A[7],
		A[6],
		A[5],
		A[4],
		A[3],
		A[2],
		A[1],
		A[0] }),
	.B({ B[7],
		B[6],
		B[5],
		B[4],
		B[3],
		B[2],
		B[1],
		B[0] }),
	.TC(1'b0),
	.PRODUCT({ N125,
		N124,
		N123,
		N122,
		N121,
		N120,
		N119,
		N118,
		N117,
		N116,
		N115,
		N114,
		N113,
		N112,
		N111,
		N110 }),
	.n135(n135),
	.n137(n137),
	.n139(n139),
	.n158(n158),
	.n157(n157),
	.n156(n156),
	.n155(n155),
	.n154(n154),
	.n153(n153),
	.n152(n152),
	.n151(n151),
	.n148(n148),
	.n149(n149),
	.n140(n140), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW_div_uns_0 (
	a, 
	b, 
	quotient, 
	remainder, 
	divide_by_0, 
	n148, 
	n158, 
	n157, 
	n140, 
	VDD, 
	VSS);
   input [7:0] a;
   input [7:0] b;
   output [7:0] quotient;
   output [7:0] remainder;
   output divide_by_0;
   input n148;
   input n158;
   input n157;
   input n140;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_RN_459_0;
   wire FE_RN_458_0;
   wire FE_RN_457_0;
   wire FE_RN_456_0;
   wire FE_RN_455_0;
   wire FE_RN_454_0;
   wire FE_RN_453_0;
   wire FE_RN_452_0;
   wire FE_RN_451_0;
   wire FE_RN_450_0;
   wire FE_RN_449_0;
   wire FE_RN_448_0;
   wire FE_RN_447_0;
   wire FE_RN_446_0;
   wire FE_RN_445_0;
   wire FE_RN_444_0;
   wire FE_RN_443_0;
   wire FE_RN_442_0;
   wire FE_RN_441_0;
   wire FE_RN_440_0;
   wire FE_RN_439_0;
   wire FE_RN_438_0;
   wire FE_RN_437_0;
   wire FE_RN_436_0;
   wire FE_RN_435_0;
   wire FE_RN_434_0;
   wire FE_RN_433_0;
   wire FE_RN_432_0;
   wire FE_RN_431_0;
   wire FE_RN_430_0;
   wire FE_RN_429_0;
   wire FE_RN_428_0;
   wire FE_RN_427_0;
   wire FE_RN_425_0;
   wire FE_RN_424_0;
   wire FE_RN_422_0;
   wire FE_RN_421_0;
   wire FE_RN_420_0;
   wire FE_RN_419_0;
   wire FE_RN_418_0;
   wire FE_RN_417_0;
   wire FE_RN_416_0;
   wire FE_RN_415_0;
   wire FE_RN_414_0;
   wire FE_RN_413_0;
   wire FE_RN_412_0;
   wire FE_RN_411_0;
   wire FE_RN_410_0;
   wire FE_RN_409_0;
   wire FE_RN_408_0;
   wire FE_RN_407_0;
   wire FE_RN_406_0;
   wire FE_RN_405_0;
   wire FE_RN_404_0;
   wire FE_RN_403_0;
   wire FE_RN_402_0;
   wire FE_RN_401_0;
   wire FE_RN_400_0;
   wire FE_RN_399_0;
   wire FE_RN_398_0;
   wire FE_RN_397_0;
   wire FE_RN_396_0;
   wire FE_RN_395_0;
   wire FE_RN_394_0;
   wire FE_RN_393_0;
   wire FE_RN_392_0;
   wire FE_RN_391_0;
   wire FE_RN_390_0;
   wire FE_RN_389_0;
   wire FE_RN_388_0;
   wire FE_RN_387_0;
   wire FE_RN_386_0;
   wire FE_RN_385_0;
   wire FE_RN_384_0;
   wire FE_RN_383_0;
   wire FE_RN_348_0;
   wire FE_RN_347_0;
   wire FE_RN_346_0;
   wire FE_RN_345_0;
   wire FE_RN_344_0;
   wire FE_RN_343_0;
   wire FE_RN_342_0;
   wire FE_RN_341_0;
   wire FE_RN_340_0;
   wire FE_RN_339_0;
   wire FE_RN_338_0;
   wire FE_RN_337_0;
   wire FE_RN_336_0;
   wire FE_RN_335_0;
   wire FE_RN_334_0;
   wire FE_RN_333_0;
   wire FE_RN_332_0;
   wire FE_RN_331_0;
   wire FE_RN_330_0;
   wire FE_RN_329_0;
   wire FE_RN_328_0;
   wire FE_RN_327_0;
   wire FE_RN_326_0;
   wire FE_RN_325_0;
   wire FE_RN_324_0;
   wire FE_RN_323_0;
   wire FE_RN_322_0;
   wire FE_RN_321_0;
   wire FE_RN_320_0;
   wire FE_RN_319_0;
   wire FE_RN_318_0;
   wire FE_RN_317_0;
   wire FE_RN_316_0;
   wire FE_RN_315_0;
   wire FE_RN_314_0;
   wire FE_RN_313_0;
   wire FE_RN_312_0;
   wire FE_RN_311_0;
   wire FE_RN_310_0;
   wire FE_RN_309_0;
   wire FE_RN_308_0;
   wire FE_RN_307_0;
   wire FE_RN_306_0;
   wire FE_RN_287_0;
   wire FE_RN_286_0;
   wire FE_RN_285_0;
   wire FE_RN_284_0;
   wire FE_RN_283_0;
   wire FE_RN_282_0;
   wire FE_RN_281_0;
   wire FE_RN_280_0;
   wire FE_RN_279_0;
   wire FE_RN_278_0;
   wire FE_RN_277_0;
   wire FE_RN_276_0;
   wire FE_RN_275_0;
   wire FE_RN_274_0;
   wire FE_RN_273_0;
   wire FE_RN_272_0;
   wire FE_RN_271_0;
   wire FE_RN_270_0;
   wire FE_RN_269_0;
   wire FE_RN_268_0;
   wire FE_RN_267_0;
   wire FE_RN_266_0;
   wire FE_RN_265_0;
   wire FE_RN_264_0;
   wire FE_RN_263_0;
   wire FE_RN_262_0;
   wire FE_RN_261_0;
   wire FE_RN_260_0;
   wire FE_RN_259_0;
   wire FE_RN_258_0;
   wire FE_RN_257_0;
   wire FE_RN_256_0;
   wire FE_RN_255_0;
   wire FE_RN_254_0;
   wire FE_RN_253_0;
   wire FE_RN_252_0;
   wire FE_RN_246_0;
   wire FE_RN_245_0;
   wire FE_RN_244_0;
   wire FE_RN_243_0;
   wire FE_RN_241_0;
   wire FE_RN_240_0;
   wire FE_RN_239_0;
   wire FE_RN_238_0;
   wire FE_RN_237_0;
   wire FE_RN_236_0;
   wire FE_RN_235_0;
   wire FE_RN_234_0;
   wire FE_RN_233_0;
   wire FE_RN_232_0;
   wire FE_RN_231_0;
   wire FE_RN_230_0;
   wire FE_RN_229_0;
   wire FE_RN_228_0;
   wire FE_RN_227_0;
   wire FE_RN_226_0;
   wire FE_RN_224_0;
   wire FE_RN_223_0;
   wire FE_RN_222_0;
   wire FE_RN_221_0;
   wire FE_RN_220_0;
   wire FE_RN_219_0;
   wire FE_RN_218_0;
   wire FE_RN_217_0;
   wire FE_RN_216_0;
   wire FE_RN_215_0;
   wire FE_RN_214_0;
   wire FE_RN_213_0;
   wire FE_RN_212_0;
   wire FE_RN_211_0;
   wire FE_RN_210_0;
   wire FE_RN_208_0;
   wire FE_RN_207_0;
   wire FE_RN_206_0;
   wire FE_RN_205_0;
   wire FE_RN_204_0;
   wire FE_RN_203_0;
   wire FE_RN_202_0;
   wire FE_RN_201_0;
   wire FE_RN_200_0;
   wire FE_RN_199_0;
   wire FE_RN_198_0;
   wire FE_RN_197_0;
   wire FE_RN_196_0;
   wire FE_RN_195_0;
   wire FE_RN_194_0;
   wire FE_RN_193_0;
   wire FE_RN_192_0;
   wire FE_RN_190_0;
   wire FE_RN_189_0;
   wire FE_RN_188_0;
   wire FE_RN_187_0;
   wire FE_RN_186_0;
   wire FE_RN_185_0;
   wire FE_RN_184_0;
   wire FE_RN_183_0;
   wire FE_RN_182_0;
   wire FE_RN_181_0;
   wire FE_RN_180_0;
   wire FE_RN_179_0;
   wire FE_RN_178_0;
   wire FE_RN_177_0;
   wire FE_RN_176_0;
   wire FE_RN_175_0;
   wire FE_RN_174_0;
   wire FE_RN_173_0;
   wire FE_RN_172_0;
   wire FE_RN_171_0;
   wire FE_RN_170_0;
   wire FE_RN_169_0;
   wire FE_RN_168_0;
   wire FE_RN_167_0;
   wire FE_RN_166_0;
   wire FE_RN_165_0;
   wire FE_RN_164_0;
   wire FE_RN_163_0;
   wire FE_RN_162_0;
   wire FE_RN_161_0;
   wire FE_RN_160_0;
   wire FE_RN_159_0;
   wire FE_RN_158_0;
   wire FE_RN_157_0;
   wire FE_RN_156_0;
   wire FE_RN_155_0;
   wire FE_RN_154_0;
   wire FE_RN_153_0;
   wire FE_RN_152_0;
   wire FE_RN_151_0;
   wire FE_RN_150_0;
   wire FE_RN_149_0;
   wire FE_RN_148_0;
   wire FE_RN_147_0;
   wire FE_RN_146_0;
   wire FE_RN_145_0;
   wire FE_RN_144_0;
   wire FE_RN_143_0;
   wire FE_RN_142_0;
   wire FE_RN_141_0;
   wire FE_RN_140_0;
   wire FE_RN_139_0;
   wire FE_RN_112_0;
   wire FE_RN_111_0;
   wire FE_RN_110_0;
   wire FE_RN_109_0;
   wire FE_RN_108_0;
   wire FE_RN_107_0;
   wire FE_RN_106_0;
   wire FE_RN_105_0;
   wire FE_RN_104_0;
   wire FE_RN_103_0;
   wire FE_RN_102_0;
   wire FE_RN_101_0;
   wire FE_RN_100_0;
   wire FE_RN_99_0;
   wire FE_RN_98_0;
   wire FE_RN_97_0;
   wire FE_RN_96_0;
   wire FE_RN_95_0;
   wire FE_RN_94_0;
   wire FE_RN_93_0;
   wire FE_RN_92_0;
   wire FE_RN_91_0;
   wire FE_RN_90_0;
   wire FE_RN_89_0;
   wire FE_RN_87_0;
   wire FE_RN_85_0;
   wire FE_RN_84_0;
   wire FE_RN_83_0;
   wire FE_RN_82_0;
   wire FE_RN_81_0;
   wire FE_RN_80_0;
   wire FE_RN_79_0;
   wire FE_RN_78_0;
   wire FE_RN_77_0;
   wire FE_RN_76_0;
   wire FE_RN_75_0;
   wire FE_RN_74_0;
   wire FE_RN_73_0;
   wire FE_RN_72_0;
   wire FE_RN_69_0;
   wire FE_RN_68_0;
   wire FE_RN_67_0;
   wire FE_RN_66_0;
   wire FE_RN_65_0;
   wire FE_RN_64_0;
   wire FE_RN_63_0;
   wire FE_RN_62_0;
   wire FE_RN_59_0;
   wire FE_RN_58_0;
   wire FE_RN_57_0;
   wire FE_RN_56_0;
   wire FE_RN_55_0;
   wire FE_RN_54_0;
   wire FE_RN_53_0;
   wire FE_RN_52_0;
   wire FE_RN_51_0;
   wire FE_RN_50_0;
   wire FE_RN_49_0;
   wire FE_RN_48_0;
   wire FE_RN_47_0;
   wire FE_RN_46_0;
   wire FE_RN_45_0;
   wire FE_RN_44_0;
   wire FE_RN_43_0;
   wire FE_RN_42_0;
   wire FE_RN_41_0;
   wire FE_RN_40_0;
   wire FE_RN_39_0;
   wire FE_RN_38_0;
   wire FE_RN_37_0;
   wire FE_RN_36_0;
   wire FE_RN_35_0;
   wire FE_RN_34_0;
   wire FE_RN_33_0;
   wire FE_RN_32_0;
   wire FE_RN_31_0;
   wire FE_RN_30_0;
   wire FE_RN_29_0;
   wire FE_RN_28_0;
   wire FE_RN_27_0;
   wire FE_RN_25_0;
   wire FE_RN_24_0;
   wire FE_RN_23_0;
   wire FE_RN_22_0;
   wire FE_RN_21_0;
   wire FE_RN_20_0;
   wire FE_RN_19_0;
   wire FE_RN_18_0;
   wire FE_RN_17_0;
   wire FE_RN_16_0;
   wire FE_RN_15_0;
   wire FE_RN_14_0;
   wire FE_RN_13_0;
   wire FE_RN_11_0;
   wire FE_RN_10_0;
   wire FE_RN_9_0;
   wire FE_RN_8_0;
   wire FE_RN_7_0;
   wire FE_RN_6_0;
   wire FE_RN_5_0;
   wire FE_RN_4_0;
   wire FE_RN_3_0;
   wire FE_RN_2_0;
   wire \u_div/SumTmp[1][0] ;
   wire \u_div/SumTmp[1][1] ;
   wire \u_div/SumTmp[1][2] ;
   wire \u_div/SumTmp[1][3] ;
   wire \u_div/SumTmp[1][4] ;
   wire \u_div/SumTmp[1][5] ;
   wire \u_div/SumTmp[1][6] ;
   wire \u_div/SumTmp[2][0] ;
   wire \u_div/SumTmp[2][1] ;
   wire \u_div/SumTmp[2][2] ;
   wire \u_div/SumTmp[2][3] ;
   wire \u_div/SumTmp[2][4] ;
   wire \u_div/SumTmp[2][5] ;
   wire \u_div/SumTmp[3][0] ;
   wire \u_div/SumTmp[3][1] ;
   wire \u_div/SumTmp[3][2] ;
   wire \u_div/SumTmp[3][3] ;
   wire \u_div/SumTmp[3][4] ;
   wire \u_div/SumTmp[4][0] ;
   wire \u_div/SumTmp[4][1] ;
   wire \u_div/SumTmp[4][2] ;
   wire \u_div/SumTmp[4][3] ;
   wire \u_div/SumTmp[5][0] ;
   wire \u_div/SumTmp[5][1] ;
   wire \u_div/SumTmp[5][2] ;
   wire \u_div/SumTmp[6][0] ;
   wire \u_div/SumTmp[6][1] ;
   wire \u_div/SumTmp[7][0] ;
   wire \u_div/CryTmp[0][1] ;
   wire \u_div/CryTmp[0][2] ;
   wire \u_div/CryTmp[0][3] ;
   wire \u_div/CryTmp[0][4] ;
   wire \u_div/CryTmp[0][5] ;
   wire \u_div/CryTmp[0][6] ;
   wire \u_div/CryTmp[0][7] ;
   wire \u_div/CryTmp[1][1] ;
   wire \u_div/CryTmp[1][6] ;
   wire \u_div/CryTmp[1][7] ;
   wire \u_div/CryTmp[2][1] ;
   wire \u_div/CryTmp[2][2] ;
   wire \u_div/CryTmp[2][3] ;
   wire \u_div/CryTmp[2][6] ;
   wire \u_div/CryTmp[3][1] ;
   wire \u_div/CryTmp[3][2] ;
   wire \u_div/CryTmp[3][3] ;
   wire \u_div/CryTmp[4][1] ;
   wire \u_div/CryTmp[4][2] ;
   wire \u_div/CryTmp[5][1] ;
   wire \u_div/CryTmp[5][2] ;
   wire \u_div/CryTmp[6][1] ;
   wire \u_div/CryTmp[7][1] ;
   wire \u_div/PartRem[1][1] ;
   wire \u_div/PartRem[1][2] ;
   wire \u_div/PartRem[1][3] ;
   wire \u_div/PartRem[1][4] ;
   wire \u_div/PartRem[1][5] ;
   wire \u_div/PartRem[1][6] ;
   wire \u_div/PartRem[1][7] ;
   wire \u_div/PartRem[2][1] ;
   wire \u_div/PartRem[2][2] ;
   wire \u_div/PartRem[2][3] ;
   wire \u_div/PartRem[2][4] ;
   wire \u_div/PartRem[2][5] ;
   wire \u_div/PartRem[2][6] ;
   wire \u_div/PartRem[3][1] ;
   wire \u_div/PartRem[3][2] ;
   wire \u_div/PartRem[3][3] ;
   wire \u_div/PartRem[3][4] ;
   wire \u_div/PartRem[3][5] ;
   wire \u_div/PartRem[4][1] ;
   wire \u_div/PartRem[4][2] ;
   wire \u_div/PartRem[4][3] ;
   wire \u_div/PartRem[4][4] ;
   wire \u_div/PartRem[5][1] ;
   wire \u_div/PartRem[5][2] ;
   wire \u_div/PartRem[5][3] ;
   wire \u_div/PartRem[6][1] ;
   wire \u_div/PartRem[6][2] ;
   wire \u_div/PartRem[7][1] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;

   // Module instantiations
   NAND2X3M FE_RC_551_0 (
	.Y(FE_RN_459_0),
	.B(FE_RN_457_0),
	.A(FE_RN_445_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_550_0 (
	.Y(FE_RN_458_0),
	.A(FE_RN_447_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_549_0 (
	.Y(FE_RN_457_0),
	.B(FE_RN_442_0),
	.A(FE_RN_458_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_548_0 (
	.Y(FE_RN_456_0),
	.C(FE_RN_457_0),
	.B(FE_RN_424_0),
	.AN(FE_RN_409_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_547_0 (
	.Y(FE_RN_455_0),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_546_0 (
	.Y(FE_RN_454_0),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_545_0 (
	.Y(FE_RN_453_0),
	.A(FE_RN_447_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_544_0 (
	.Y(FE_RN_452_0),
	.B0(FE_RN_453_0),
	.A1N(FE_RN_454_0),
	.A0N(FE_RN_455_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_543_0 (
	.Y(FE_RN_451_0),
	.A(FE_RN_452_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_542_0 (
	.Y(FE_RN_450_0),
	.B(FE_RN_415_0),
	.A(FE_RN_409_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_541_0 (
	.Y(FE_RN_449_0),
	.B(FE_RN_424_0),
	.A(FE_RN_450_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_540_0 (
	.Y(FE_RN_448_0),
	.C(FE_RN_427_0),
	.B(FE_RN_451_0),
	.A(FE_RN_449_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_539_0 (
	.Y(\u_div/SumTmp[1][5] ),
	.C(FE_RN_459_0),
	.B(FE_RN_456_0),
	.A(FE_RN_448_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKAND2X4M FE_RC_538_0 (
	.Y(FE_RN_447_0),
	.B(n13),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_537_0 (
	.Y(FE_RN_446_0),
	.A(FE_RN_447_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X4M FE_RC_536_0 (
	.Y(FE_RN_445_0),
	.B0(FE_RN_427_0),
	.A1N(FE_RN_424_0),
	.A0(FE_RN_415_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_535_0 (
	.Y(FE_RN_444_0),
	.B(FE_RN_442_0),
	.A(FE_RN_445_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_534_0 (
	.Y(FE_RN_443_0),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_533_0 (
	.Y(FE_RN_442_0),
	.B(FE_RN_443_0),
	.AN(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_532_0 (
	.Y(FE_RN_441_0),
	.C(FE_RN_442_0),
	.B(FE_RN_424_0),
	.AN(FE_RN_409_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_531_0 (
	.Y(\u_div/CryTmp[1][6] ),
	.C(FE_RN_446_0),
	.B(FE_RN_444_0),
	.A(FE_RN_441_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_530_0 (
	.Y(FE_RN_440_0),
	.A(FE_RN_415_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_529_0 (
	.Y(FE_RN_439_0),
	.B(FE_RN_440_0),
	.A(FE_RN_436_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_528_0 (
	.Y(FE_RN_438_0),
	.A(FE_RN_409_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_527_0 (
	.Y(FE_RN_437_0),
	.A(FE_RN_428_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_526_0 (
	.Y(FE_RN_436_0),
	.B(FE_RN_424_0),
	.A(FE_RN_437_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_525_0 (
	.Y(FE_RN_435_0),
	.B(FE_RN_438_0),
	.A(FE_RN_436_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_524_0 (
	.Y(FE_RN_434_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_523_0 (
	.Y(FE_RN_433_0),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_522_0 (
	.Y(FE_RN_432_0),
	.A(FE_RN_428_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_521_0 (
	.Y(FE_RN_431_0),
	.B0(FE_RN_432_0),
	.A1N(FE_RN_433_0),
	.A0N(FE_RN_434_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_520_0 (
	.Y(FE_RN_430_0),
	.A(FE_RN_431_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_519_0 (
	.Y(FE_RN_429_0),
	.C(FE_RN_415_0),
	.B(FE_RN_409_0),
	.A(FE_RN_430_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_518_0 (
	.Y(\u_div/SumTmp[1][4] ),
	.C(FE_RN_439_0),
	.B(FE_RN_435_0),
	.A(FE_RN_429_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKAND2X4M FE_RC_517_0 (
	.Y(FE_RN_428_0),
	.B(n14),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_516_0 (
	.Y(FE_RN_427_0),
	.A(FE_RN_428_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_514_0 (
	.Y(FE_RN_425_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_513_0 (
	.Y(FE_RN_424_0),
	.B(FE_RN_425_0),
	.AN(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_510_0 (
	.Y(FE_RN_422_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_509_0 (
	.Y(FE_RN_421_0),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_508_0 (
	.Y(FE_RN_420_0),
	.A(FE_RN_416_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_507_0 (
	.Y(FE_RN_419_0),
	.B0(FE_RN_420_0),
	.A1N(FE_RN_421_0),
	.A0N(FE_RN_422_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_506_0 (
	.Y(FE_RN_418_0),
	.A(FE_RN_413_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_505_0 (
	.Y(FE_RN_417_0),
	.B(FE_RN_418_0),
	.A(FE_RN_416_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_504_0 (
	.Y(\u_div/SumTmp[1][3] ),
	.S0(FE_RN_410_0),
	.B(FE_RN_417_0),
	.A(FE_RN_419_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKAND2X6M FE_RC_503_0 (
	.Y(FE_RN_416_0),
	.B(n15),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_502_0 (
	.Y(FE_RN_415_0),
	.A(FE_RN_416_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_501_0 (
	.Y(FE_RN_414_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_500_0 (
	.Y(FE_RN_413_0),
	.B(FE_RN_414_0),
	.AN(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_499_0 (
	.Y(FE_RN_412_0),
	.A(FE_RN_393_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_498_0 (
	.Y(FE_RN_411_0),
	.B(\u_div/PartRem[2][2] ),
	.A(FE_RN_412_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_497_0 (
	.Y(FE_RN_410_0),
	.B(FE_RN_383_0),
	.A(FE_RN_411_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_496_0 (
	.Y(FE_RN_409_0),
	.B(FE_RN_413_0),
	.A(FE_RN_410_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX6M FE_RC_494_0 (
	.Y(quotient[2]),
	.A(FE_RN_389_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_493_0 (
	.Y(FE_RN_408_0),
	.A(\u_div/SumTmp[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_492_0 (
	.Y(FE_RN_407_0),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_491_0 (
	.Y(\u_div/PartRem[2][1] ),
	.S0(FE_RN_389_0),
	.B(FE_RN_407_0),
	.A(FE_RN_408_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_490_0 (
	.Y(FE_RN_406_0),
	.A(FE_RN_384_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_489_0 (
	.Y(FE_RN_405_0),
	.A(\u_div/CryTmp[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_488_0 (
	.Y(FE_RN_404_0),
	.A(FE_RN_386_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M FE_RC_487_0 (
	.Y(FE_RN_403_0),
	.B0(FE_RN_404_0),
	.A1(FE_RN_405_0),
	.A0(FE_RN_392_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X4M FE_RC_486_0 (
	.Y(FE_RN_402_0),
	.B(n16),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_485_0 (
	.Y(\u_div/SumTmp[1][2] ),
	.S0(FE_RN_402_0),
	.B(FE_RN_403_0),
	.A(FE_RN_406_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_484_0 (
	.Y(FE_RN_401_0),
	.A(\u_div/CryTmp[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X8M FE_RC_483_0 (
	.Y(FE_RN_400_0),
	.B(n17),
	.A(FE_RN_388_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_482_0 (
	.Y(FE_RN_399_0),
	.B(FE_RN_401_0),
	.A(FE_RN_400_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_481_0 (
	.Y(FE_RN_398_0),
	.B(FE_RN_392_0),
	.A(FE_RN_386_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_480_0 (
	.Y(FE_RN_397_0),
	.B(\u_div/CryTmp[1][1] ),
	.A(FE_RN_398_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_479_0 (
	.Y(\u_div/SumTmp[1][1] ),
	.B(FE_RN_399_0),
	.A(FE_RN_397_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_478_0 (
	.Y(FE_RN_396_0),
	.A(\u_div/CryTmp[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_477_0 (
	.Y(FE_RN_395_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_476_0 (
	.Y(FE_RN_394_0),
	.B(FE_RN_395_0),
	.A(FE_RN_392_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X8M FE_RC_475_0 (
	.Y(FE_RN_393_0),
	.B0(FE_RN_394_0),
	.A1N(FE_RN_396_0),
	.A0(FE_RN_386_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X6M FE_RC_474_0 (
	.Y(FE_RN_392_0),
	.B(n17),
	.A(FE_RN_388_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_473_0 (
	.Y(FE_RN_391_0),
	.A(\u_div/SumTmp[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_472_0 (
	.Y(FE_RN_390_0),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X8M FE_RC_471_0 (
	.Y(FE_RN_389_0),
	.B(n21),
	.A(\u_div/CryTmp[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X6M FE_RC_470_0 (
	.Y(FE_RN_388_0),
	.S0(FE_RN_389_0),
	.B(FE_RN_390_0),
	.A(FE_RN_391_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_469_0 (
	.Y(FE_RN_387_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_468_0 (
	.Y(FE_RN_386_0),
	.B(FE_RN_387_0),
	.AN(FE_RN_388_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X8M FE_RC_467_0 (
	.Y(FE_RN_385_0),
	.B(\u_div/CryTmp[1][1] ),
	.A(FE_RN_386_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_466_0 (
	.Y(FE_RN_384_0),
	.B(FE_RN_392_0),
	.A(FE_RN_385_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_465_0 (
	.Y(FE_RN_383_0),
	.B(n16),
	.A(FE_RN_384_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X6M FE_RC_422_0 (
	.Y(\u_div/CryTmp[2][3] ),
	.B(FE_RN_269_0),
	.A(FE_RN_276_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_421_0 (
	.Y(FE_RN_348_0),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_420_0 (
	.Y(FE_RN_347_0),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_419_0 (
	.Y(FE_RN_346_0),
	.A(FE_RN_341_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_418_0 (
	.Y(FE_RN_345_0),
	.B0(FE_RN_346_0),
	.A1N(FE_RN_347_0),
	.A0N(FE_RN_348_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_417_0 (
	.Y(FE_RN_344_0),
	.A(FE_RN_338_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_416_0 (
	.Y(FE_RN_343_0),
	.B(FE_RN_344_0),
	.A(FE_RN_341_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_415_0 (
	.Y(\u_div/SumTmp[2][5] ),
	.S0(FE_RN_332_0),
	.B(FE_RN_343_0),
	.A(FE_RN_345_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_414_0 (
	.Y(FE_RN_342_0),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_413_0 (
	.Y(FE_RN_341_0),
	.B(FE_RN_342_0),
	.AN(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_412_0 (
	.Y(FE_RN_340_0),
	.A(FE_RN_341_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_411_0 (
	.Y(FE_RN_339_0),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_410_0 (
	.Y(FE_RN_338_0),
	.B(FE_RN_339_0),
	.AN(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_409_0 (
	.Y(FE_RN_337_0),
	.B(FE_RN_276_0),
	.A(FE_RN_269_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_408_0 (
	.Y(FE_RN_336_0),
	.C(FE_RN_337_0),
	.B(FE_RN_309_0),
	.A(FE_RN_306_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_407_0 (
	.Y(FE_RN_335_0),
	.A(FE_RN_315_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_406_0 (
	.Y(FE_RN_334_0),
	.A(FE_RN_312_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X3M FE_RC_405_0 (
	.Y(FE_RN_333_0),
	.B(FE_RN_335_0),
	.A(FE_RN_334_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_404_0 (
	.Y(FE_RN_332_0),
	.B(FE_RN_336_0),
	.A(FE_RN_333_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_403_0 (
	.Y(FE_RN_331_0),
	.B(FE_RN_338_0),
	.A(FE_RN_332_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_402_0 (
	.Y(\u_div/CryTmp[2][6] ),
	.B(FE_RN_340_0),
	.A(FE_RN_331_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_401_0 (
	.Y(FE_RN_330_0),
	.A(FE_RN_314_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_400_0 (
	.Y(FE_RN_329_0),
	.B(FE_RN_330_0),
	.A(FE_RN_322_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_399_0 (
	.Y(FE_RN_328_0),
	.B(n14),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_398_0 (
	.Y(FE_RN_327_0),
	.A(\u_div/CryTmp[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_397_0 (
	.Y(FE_RN_326_0),
	.B(FE_RN_327_0),
	.A(FE_RN_314_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_396_0 (
	.Y(FE_RN_325_0),
	.B(FE_RN_306_0),
	.A(FE_RN_326_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_395_0 (
	.Y(FE_RN_324_0),
	.B(FE_RN_328_0),
	.A(FE_RN_325_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_394_0 (
	.Y(FE_RN_323_0),
	.B(n14),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_393_0 (
	.Y(FE_RN_322_0),
	.B(FE_RN_323_0),
	.A(FE_RN_309_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_392_0 (
	.Y(FE_RN_321_0),
	.C(\u_div/CryTmp[2][3] ),
	.B(FE_RN_306_0),
	.A(FE_RN_322_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_391_0 (
	.Y(\u_div/SumTmp[2][4] ),
	.C(FE_RN_329_0),
	.B(FE_RN_324_0),
	.A(FE_RN_321_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_390_0 (
	.Y(FE_RN_320_0),
	.B(n15),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_389_0 (
	.Y(FE_RN_319_0),
	.A(\u_div/CryTmp[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_388_0 (
	.Y(FE_RN_318_0),
	.B(FE_RN_319_0),
	.AN(FE_RN_320_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_387_0 (
	.Y(FE_RN_317_0),
	.B(FE_RN_314_0),
	.A(FE_RN_306_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_386_0 (
	.Y(FE_RN_316_0),
	.B(\u_div/CryTmp[2][3] ),
	.A(FE_RN_317_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_385_0 (
	.Y(\u_div/SumTmp[2][3] ),
	.B(FE_RN_318_0),
	.A(FE_RN_316_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_384_0 (
	.Y(FE_RN_315_0),
	.B(n14),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_383_0 (
	.Y(FE_RN_314_0),
	.B(n15),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_382_0 (
	.Y(FE_RN_313_0),
	.A(FE_RN_314_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_381_0 (
	.Y(FE_RN_312_0),
	.B(FE_RN_313_0),
	.A(FE_RN_309_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_380_0 (
	.Y(FE_RN_311_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_379_0 (
	.Y(FE_RN_310_0),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_378_0 (
	.Y(FE_RN_309_0),
	.B(FE_RN_311_0),
	.A(FE_RN_310_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_377_0 (
	.Y(FE_RN_308_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_376_0 (
	.Y(FE_RN_307_0),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_375_0 (
	.Y(FE_RN_306_0),
	.B(FE_RN_308_0),
	.A(FE_RN_307_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_353_0 (
	.Y(quotient[3]),
	.B(FE_RN_244_0),
	.A(FE_RN_258_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_352_0 (
	.Y(FE_RN_287_0),
	.A(FE_RN_271_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_351_0 (
	.Y(FE_RN_286_0),
	.A(FE_RN_274_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_350_0 (
	.Y(\u_div/PartRem[3][2] ),
	.B(FE_RN_287_0),
	.A(FE_RN_286_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_349_0 (
	.Y(FE_RN_285_0),
	.A(FE_RN_279_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_348_0 (
	.Y(FE_RN_284_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M FE_RC_347_0 (
	.Y(FE_RN_283_0),
	.B1(\u_div/SumTmp[3][1] ),
	.B0(FE_RN_284_0),
	.A1N(\u_div/SumTmp[3][1] ),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_346_0 (
	.Y(FE_RN_282_0),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_345_0 (
	.Y(FE_RN_281_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M FE_RC_344_0 (
	.Y(FE_RN_280_0),
	.B1(\u_div/PartRem[4][1] ),
	.B0(FE_RN_281_0),
	.A1(n16),
	.A0(FE_RN_282_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X4M FE_RC_343_0 (
	.Y(FE_RN_279_0),
	.B1(FE_RN_280_0),
	.B0(FE_RN_272_0),
	.A1N(FE_RN_272_0),
	.A0N(FE_RN_283_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_342_0 (
	.Y(FE_RN_278_0),
	.A(FE_RN_279_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_341_0 (
	.Y(FE_RN_277_0),
	.B(\u_div/CryTmp[2][2] ),
	.A(FE_RN_278_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_340_0 (
	.Y(\u_div/SumTmp[2][2] ),
	.B0(FE_RN_277_0),
	.A1(\u_div/CryTmp[2][2] ),
	.A0(FE_RN_285_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X6M FE_RC_339_0 (
	.Y(FE_RN_276_0),
	.B0(n16),
	.A1(FE_RN_271_0),
	.A0(FE_RN_274_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_338_0 (
	.Y(FE_RN_275_0),
	.A(\u_div/PartRem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_337_0 (
	.Y(FE_RN_274_0),
	.B(FE_RN_275_0),
	.A(FE_RN_272_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_336_0 (
	.Y(FE_RN_273_0),
	.A(FE_RN_274_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_335_0 (
	.Y(FE_RN_272_0),
	.B(FE_RN_258_0),
	.A(FE_RN_244_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_334_0 (
	.Y(FE_RN_271_0),
	.B(\u_div/SumTmp[3][1] ),
	.A(FE_RN_272_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_333_0 (
	.Y(FE_RN_270_0),
	.B(n16),
	.A(FE_RN_271_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X4M FE_RC_332_0 (
	.Y(FE_RN_269_0),
	.B0(\u_div/CryTmp[2][2] ),
	.A1N(FE_RN_270_0),
	.A0N(FE_RN_273_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_329_0 (
	.Y(FE_RN_268_0),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_328_0 (
	.Y(FE_RN_267_0),
	.A(\u_div/SumTmp[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_327_0 (
	.Y(\u_div/PartRem[3][1] ),
	.S0(FE_RN_257_0),
	.B(FE_RN_267_0),
	.A(FE_RN_268_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2X8M FE_RC_326_0 (
	.Y(FE_RN_266_0),
	.B1(FE_RN_263_0),
	.B0(a[3]),
	.A1N(a[3]),
	.A0N(FE_RN_263_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_325_0 (
	.Y(FE_RN_265_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_324_0 (
	.Y(FE_RN_264_0),
	.A(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X8M FE_RC_323_0 (
	.Y(FE_RN_263_0),
	.B0(FE_RN_254_0),
	.A1(FE_RN_264_0),
	.A0(FE_RN_265_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_322_0 (
	.Y(FE_RN_262_0),
	.B(\u_div/SumTmp[3][0] ),
	.A(FE_RN_263_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_321_0 (
	.Y(FE_RN_261_0),
	.B0(FE_RN_262_0),
	.A1(\u_div/SumTmp[3][0] ),
	.A0(FE_RN_263_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_320_0 (
	.Y(\u_div/SumTmp[2][1] ),
	.S0(FE_RN_257_0),
	.B(FE_RN_261_0),
	.A(FE_RN_266_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_319_0 (
	.Y(FE_RN_260_0),
	.A(FE_RN_243_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX4M FE_RC_318_0 (
	.Y(FE_RN_259_0),
	.B(FE_RN_260_0),
	.AN(FE_RN_230_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_317_0 (
	.Y(FE_RN_258_0),
	.B(FE_RN_226_0),
	.A(FE_RN_259_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X12M FE_RC_316_0 (
	.Y(FE_RN_257_0),
	.B(FE_RN_244_0),
	.A(FE_RN_258_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_315_0 (
	.Y(FE_RN_256_0),
	.S0(FE_RN_257_0),
	.B(\u_div/SumTmp[3][0] ),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_314_0 (
	.Y(FE_RN_255_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_313_0 (
	.Y(FE_RN_254_0),
	.B(FE_RN_255_0),
	.AN(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_312_0 (
	.Y(FE_RN_253_0),
	.A(\u_div/CryTmp[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_311_0 (
	.Y(FE_RN_252_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X8M FE_RC_310_0 (
	.Y(\u_div/CryTmp[2][2] ),
	.B1(FE_RN_252_0),
	.B0(FE_RN_253_0),
	.A1N(FE_RN_254_0),
	.A0(FE_RN_256_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_302_0 (
	.Y(FE_RN_246_0),
	.B(n13),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_301_0 (
	.Y(FE_RN_245_0),
	.A(FE_RN_233_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X5M FE_RC_300_0 (
	.Y(FE_RN_244_0),
	.B(FE_RN_246_0),
	.A(FE_RN_245_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_299_0 (
	.Y(FE_RN_243_0),
	.B(n13),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_296_0 (
	.Y(\u_div/CryTmp[3][3] ),
	.B(FE_RN_229_0),
	.A(FE_RN_199_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_295_0 (
	.Y(FE_RN_241_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_294_0 (
	.Y(FE_RN_240_0),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_293_0 (
	.Y(FE_RN_239_0),
	.A(FE_RN_234_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_292_0 (
	.Y(FE_RN_238_0),
	.B0(FE_RN_239_0),
	.A1N(FE_RN_240_0),
	.A0N(FE_RN_241_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_291_0 (
	.Y(FE_RN_237_0),
	.A(FE_RN_230_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_290_0 (
	.Y(FE_RN_236_0),
	.B(FE_RN_237_0),
	.A(FE_RN_234_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_289_0 (
	.Y(\u_div/SumTmp[3][4] ),
	.S0(FE_RN_226_0),
	.B(FE_RN_236_0),
	.A(FE_RN_238_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_288_0 (
	.Y(FE_RN_235_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_287_0 (
	.Y(FE_RN_234_0),
	.B(FE_RN_235_0),
	.AN(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_286_0 (
	.Y(FE_RN_233_0),
	.A(FE_RN_234_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_285_0 (
	.Y(FE_RN_232_0),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M FE_RC_284_0 (
	.Y(FE_RN_231_0),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_283_0 (
	.Y(FE_RN_230_0),
	.B(FE_RN_232_0),
	.A(FE_RN_231_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_282_0 (
	.Y(FE_RN_229_0),
	.B(\u_div/CryTmp[3][2] ),
	.A(FE_RN_192_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_281_0 (
	.Y(FE_RN_228_0),
	.B(FE_RN_199_0),
	.A(FE_RN_229_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_280_0 (
	.Y(FE_RN_227_0),
	.B(FE_RN_210_0),
	.A(FE_RN_228_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_279_0 (
	.Y(FE_RN_226_0),
	.B(FE_RN_215_0),
	.A(FE_RN_227_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_276_0 (
	.Y(FE_RN_224_0),
	.A(FE_RN_212_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_275_0 (
	.Y(FE_RN_223_0),
	.A(FE_RN_214_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_274_0 (
	.Y(\u_div/PartRem[4][3] ),
	.B(FE_RN_224_0),
	.A(FE_RN_223_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_273_0 (
	.Y(FE_RN_222_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_272_0 (
	.Y(FE_RN_221_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_271_0 (
	.Y(FE_RN_220_0),
	.B1(FE_RN_221_0),
	.B0(\u_div/SumTmp[4][2] ),
	.A1N(\u_div/SumTmp[4][2] ),
	.A0N(FE_RN_222_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_270_0 (
	.Y(FE_RN_219_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_269_0 (
	.Y(FE_RN_218_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_268_0 (
	.Y(FE_RN_217_0),
	.B1(FE_RN_218_0),
	.B0(\u_div/PartRem[5][2] ),
	.A1N(\u_div/PartRem[5][2] ),
	.A0N(FE_RN_219_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M FE_RC_267_0 (
	.Y(FE_RN_216_0),
	.B1(FE_RN_217_0),
	.B0(quotient[4]),
	.A1N(quotient[4]),
	.A0(FE_RN_220_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X4M FE_RC_266_0 (
	.Y(\u_div/SumTmp[3][3] ),
	.B1(\u_div/CryTmp[3][3] ),
	.B0(FE_RN_216_0),
	.A1N(FE_RN_216_0),
	.A0N(\u_div/CryTmp[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_265_0 (
	.Y(FE_RN_215_0),
	.B0(n15),
	.A1(FE_RN_214_0),
	.A0(FE_RN_212_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M FE_RC_264_0 (
	.Y(FE_RN_214_0),
	.B(quotient[4]),
	.A(\u_div/SumTmp[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_263_0 (
	.Y(FE_RN_213_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M FE_RC_262_0 (
	.Y(FE_RN_212_0),
	.B(quotient[4]),
	.AN(\u_div/PartRem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_261_0 (
	.Y(FE_RN_211_0),
	.A(FE_RN_212_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_260_0 (
	.Y(FE_RN_210_0),
	.C(FE_RN_211_0),
	.B(FE_RN_213_0),
	.AN(FE_RN_214_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_257_0 (
	.Y(FE_RN_208_0),
	.A(FE_RN_194_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_256_0 (
	.Y(\u_div/PartRem[4][2] ),
	.B(FE_RN_208_0),
	.AN(FE_RN_197_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_255_0 (
	.Y(FE_RN_207_0),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_254_0 (
	.Y(FE_RN_206_0),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_253_0 (
	.Y(FE_RN_205_0),
	.B1(n16),
	.B0(FE_RN_206_0),
	.A1N(FE_RN_207_0),
	.A0N(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_252_0 (
	.Y(FE_RN_204_0),
	.A(\u_div/SumTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_251_0 (
	.Y(FE_RN_203_0),
	.A(\u_div/SumTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_250_0 (
	.Y(FE_RN_202_0),
	.B1(n16),
	.B0(FE_RN_203_0),
	.A1N(FE_RN_204_0),
	.A0N(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X6M FE_RC_249_0 (
	.Y(FE_RN_201_0),
	.S0(quotient[4]),
	.B(FE_RN_202_0),
	.A(FE_RN_205_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_248_0 (
	.Y(FE_RN_200_0),
	.B(\u_div/CryTmp[3][2] ),
	.A(FE_RN_201_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_247_0 (
	.Y(\u_div/SumTmp[3][2] ),
	.B0(FE_RN_200_0),
	.A1(\u_div/CryTmp[3][2] ),
	.A0(FE_RN_201_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X8M FE_RC_246_0 (
	.Y(FE_RN_199_0),
	.B0(n16),
	.A1(FE_RN_194_0),
	.A0(FE_RN_197_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_245_0 (
	.Y(FE_RN_198_0),
	.A(\u_div/PartRem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X8M FE_RC_244_0 (
	.Y(FE_RN_197_0),
	.B(quotient[4]),
	.A(FE_RN_198_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_243_0 (
	.Y(FE_RN_196_0),
	.A(FE_RN_197_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_242_0 (
	.Y(FE_RN_195_0),
	.A(\u_div/SumTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_241_0 (
	.Y(FE_RN_194_0),
	.B(FE_RN_195_0),
	.AN(quotient[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_240_0 (
	.Y(FE_RN_193_0),
	.B(n16),
	.A(FE_RN_194_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_239_0 (
	.Y(FE_RN_192_0),
	.B(FE_RN_196_0),
	.A(FE_RN_193_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_236_0 (
	.Y(\u_div/PartRem[4][1] ),
	.S0(FE_RN_165_0),
	.B(FE_RN_168_0),
	.A(FE_RN_169_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_235_0 (
	.Y(FE_RN_190_0),
	.A(\u_div/CryTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_234_0 (
	.Y(FE_RN_189_0),
	.A(\u_div/CryTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X8M FE_RC_233_0 (
	.Y(FE_RN_188_0),
	.B1(n17),
	.B0(FE_RN_169_0),
	.A1N(FE_RN_169_0),
	.A0N(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_232_0 (
	.Y(FE_RN_187_0),
	.B(FE_RN_189_0),
	.A(FE_RN_188_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_231_0 (
	.Y(FE_RN_186_0),
	.B0(FE_RN_187_0),
	.A1(FE_RN_190_0),
	.A0(FE_RN_188_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_230_0 (
	.Y(FE_RN_185_0),
	.A(FE_RN_171_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_229_0 (
	.Y(FE_RN_184_0),
	.B0(FE_RN_185_0),
	.A1(\u_div/CryTmp[3][1] ),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_228_0 (
	.Y(FE_RN_183_0),
	.A(FE_RN_176_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_227_0 (
	.Y(FE_RN_182_0),
	.B(FE_RN_183_0),
	.A(FE_RN_171_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_226_0 (
	.Y(FE_RN_181_0),
	.A(FE_RN_168_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X3M FE_RC_225_0 (
	.Y(FE_RN_180_0),
	.S0(FE_RN_181_0),
	.B(FE_RN_182_0),
	.A(FE_RN_184_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_224_0 (
	.Y(FE_RN_179_0),
	.B(FE_RN_165_0),
	.A(FE_RN_180_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X4M FE_RC_223_0 (
	.Y(\u_div/SumTmp[3][1] ),
	.B0(FE_RN_179_0),
	.A1N(FE_RN_186_0),
	.A0(FE_RN_165_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_222_0 (
	.Y(FE_RN_178_0),
	.B(FE_RN_169_0),
	.AN(FE_RN_176_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_221_0 (
	.Y(FE_RN_177_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_220_0 (
	.Y(FE_RN_176_0),
	.B(FE_RN_177_0),
	.AN(\u_div/CryTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_219_0 (
	.Y(FE_RN_175_0),
	.A(FE_RN_176_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_218_0 (
	.Y(FE_RN_174_0),
	.B(FE_RN_168_0),
	.A(FE_RN_175_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_217_0 (
	.Y(FE_RN_173_0),
	.B(FE_RN_165_0),
	.A(FE_RN_174_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_216_0 (
	.Y(FE_RN_172_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_215_0 (
	.Y(FE_RN_171_0),
	.B(FE_RN_172_0),
	.AN(\u_div/CryTmp[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_214_0 (
	.Y(FE_RN_170_0),
	.A(FE_RN_171_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X4M FE_RC_213_0 (
	.Y(\u_div/CryTmp[3][2] ),
	.C0(FE_RN_170_0),
	.B0(FE_RN_173_0),
	.A1N(FE_RN_178_0),
	.A0(FE_RN_165_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X6M FE_RC_212_0 (
	.Y(quotient[4]),
	.B(FE_RN_166_0),
	.A(FE_RN_160_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_211_0 (
	.Y(FE_RN_169_0),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_210_0 (
	.Y(FE_RN_168_0),
	.A(\u_div/SumTmp[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_209_0 (
	.Y(FE_RN_167_0),
	.A(FE_RN_162_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_208_0 (
	.Y(FE_RN_166_0),
	.B(FE_RN_167_0),
	.AN(FE_RN_163_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_207_0 (
	.Y(FE_RN_165_0),
	.B(FE_RN_160_0),
	.A(FE_RN_166_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_205_0 (
	.Y(FE_RN_164_0),
	.A(FE_RN_140_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X4M FE_RC_204_0 (
	.Y(FE_RN_163_0),
	.B1(FE_RN_164_0),
	.B0(n15),
	.A1(\u_div/PartRem[5][3] ),
	.A0(FE_RN_139_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_203_0 (
	.Y(FE_RN_162_0),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_202_0 (
	.Y(FE_RN_161_0),
	.A(FE_RN_144_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_201_0 (
	.Y(FE_RN_160_0),
	.B(n20),
	.A(FE_RN_161_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_199_0 (
	.Y(FE_RN_159_0),
	.A(\u_div/PartRem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M FE_RC_198_0 (
	.Y(\u_div/PartRem[5][2] ),
	.B1(quotient[5]),
	.B0(FE_RN_159_0),
	.A1N(\u_div/SumTmp[5][1] ),
	.A0N(quotient[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_197_0 (
	.Y(FE_RN_158_0),
	.A(FE_RN_140_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_196_0 (
	.Y(FE_RN_157_0),
	.B0(FE_RN_158_0),
	.A1(\u_div/CryTmp[4][2] ),
	.A0(FE_RN_145_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_195_0 (
	.Y(FE_RN_156_0),
	.A(\u_div/CryTmp[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_194_0 (
	.Y(FE_RN_155_0),
	.A(FE_RN_145_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_193_0 (
	.Y(FE_RN_154_0),
	.B0(FE_RN_155_0),
	.A1(FE_RN_156_0),
	.A0(FE_RN_140_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_192_0 (
	.Y(FE_RN_153_0),
	.B(n15),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_191_0 (
	.Y(FE_RN_152_0),
	.B(FE_RN_153_0),
	.AN(FE_RN_154_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_190_0 (
	.Y(\u_div/SumTmp[4][3] ),
	.B0(FE_RN_152_0),
	.A1(FE_RN_153_0),
	.A0(FE_RN_157_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_189_0 (
	.Y(FE_RN_151_0),
	.B(n16),
	.A(FE_RN_141_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M FE_RC_188_0 (
	.Y(FE_RN_150_0),
	.B0(FE_RN_151_0),
	.A1(n16),
	.A0(FE_RN_141_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_187_0 (
	.Y(FE_RN_149_0),
	.B(FE_RN_140_0),
	.A(FE_RN_145_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_186_0 (
	.Y(FE_RN_148_0),
	.B(\u_div/CryTmp[4][2] ),
	.A(FE_RN_149_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X3M FE_RC_185_0 (
	.Y(\u_div/SumTmp[4][2] ),
	.B0(FE_RN_148_0),
	.A1(\u_div/CryTmp[4][2] ),
	.A0(FE_RN_150_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X3M FE_RC_184_0 (
	.Y(FE_RN_147_0),
	.B(n15),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_183_0 (
	.Y(FE_RN_146_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_182_0 (
	.Y(FE_RN_145_0),
	.B(FE_RN_146_0),
	.AN(FE_RN_141_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_181_0 (
	.Y(FE_RN_144_0),
	.C(\u_div/CryTmp[4][2] ),
	.B(FE_RN_145_0),
	.AN(FE_RN_147_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_180_0 (
	.Y(FE_RN_143_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_179_0 (
	.Y(FE_RN_142_0),
	.B(quotient[5]),
	.A(\u_div/SumTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X4M FE_RC_178_0 (
	.Y(FE_RN_141_0),
	.B0(FE_RN_142_0),
	.A1N(\u_div/PartRem[6][1] ),
	.A0(quotient[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X6M FE_RC_177_0 (
	.Y(FE_RN_140_0),
	.B(n16),
	.A(FE_RN_141_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_176_0 (
	.Y(FE_RN_139_0),
	.B(FE_RN_143_0),
	.A(FE_RN_140_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_143_0 (
	.Y(FE_RN_112_0),
	.A(FE_RN_99_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX4M FE_RC_142_0 (
	.Y(\u_div/PartRem[5][1] ),
	.D(FE_RN_93_0),
	.C(FE_RN_85_0),
	.B(FE_RN_75_0),
	.AN(FE_RN_112_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_141_0 (
	.Y(FE_RN_111_0),
	.A(FE_RN_99_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX4M FE_RC_140_0 (
	.Y(FE_RN_110_0),
	.D(FE_RN_93_0),
	.C(FE_RN_85_0),
	.B(FE_RN_75_0),
	.AN(FE_RN_111_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_139_0 (
	.Y(FE_RN_109_0),
	.B(FE_RN_106_0),
	.A(FE_RN_110_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_138_0 (
	.Y(FE_RN_108_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_137_0 (
	.Y(FE_RN_107_0),
	.A(\u_div/CryTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_136_0 (
	.Y(FE_RN_106_0),
	.B0(FE_RN_95_0),
	.A1(FE_RN_107_0),
	.A0(FE_RN_108_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_135_0 (
	.Y(FE_RN_105_0),
	.A(FE_RN_106_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_134_0 (
	.Y(FE_RN_104_0),
	.A(FE_RN_92_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_133_0 (
	.Y(FE_RN_103_0),
	.C(FE_RN_105_0),
	.B(FE_RN_99_0),
	.A(FE_RN_104_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_132_0 (
	.Y(\u_div/SumTmp[4][1] ),
	.B(FE_RN_109_0),
	.A(FE_RN_103_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_131_0 (
	.Y(FE_RN_102_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_130_0 (
	.Y(FE_RN_101_0),
	.B(FE_RN_102_0),
	.A(FE_RN_99_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_129_0 (
	.Y(FE_RN_100_0),
	.B(\u_div/CryTmp[4][1] ),
	.A(FE_RN_101_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X5M FE_RC_128_0 (
	.Y(FE_RN_99_0),
	.B(a[5]),
	.A(FE_RN_69_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_127_0 (
	.Y(FE_RN_98_0),
	.A(FE_RN_99_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_126_0 (
	.Y(FE_RN_97_0),
	.B(n17),
	.A(FE_RN_98_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_125_0 (
	.Y(FE_RN_96_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX4M FE_RC_124_0 (
	.Y(FE_RN_95_0),
	.B(FE_RN_96_0),
	.AN(\u_div/CryTmp[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX8M FE_RC_123_0 (
	.Y(FE_RN_94_0),
	.B(FE_RN_89_0),
	.AN(FE_RN_87_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_122_0 (
	.Y(FE_RN_93_0),
	.B(FE_RN_94_0),
	.AN(FE_RN_55_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_121_0 (
	.Y(FE_RN_92_0),
	.C(FE_RN_75_0),
	.B(FE_RN_85_0),
	.A(FE_RN_93_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_120_0 (
	.Y(FE_RN_91_0),
	.B(FE_RN_95_0),
	.A(FE_RN_92_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_119_0 (
	.Y(\u_div/CryTmp[4][2] ),
	.C(FE_RN_100_0),
	.B(FE_RN_97_0),
	.A(FE_RN_91_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_118_0 (
	.Y(FE_RN_90_0),
	.A(FE_RN_69_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X8M FE_RC_117_0 (
	.Y(quotient[5]),
	.B1(FE_RN_55_0),
	.B0(FE_RN_69_0),
	.A1N(FE_RN_90_0),
	.A0(FE_RN_77_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_116_0 (
	.Y(FE_RN_89_0),
	.A(\u_div/SumTmp[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_114_0 (
	.Y(FE_RN_87_0),
	.A(FE_RN_69_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_112_0 (
	.Y(FE_RN_85_0),
	.C(FE_RN_55_0),
	.B(a[5]),
	.A(FE_RN_77_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_111_0 (
	.Y(FE_RN_84_0),
	.A(FE_RN_69_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_110_0 (
	.Y(FE_RN_83_0),
	.A(FE_RN_72_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M FE_RC_109_0 (
	.Y(FE_RN_82_0),
	.B(FE_RN_83_0),
	.AN(FE_RN_73_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_108_0 (
	.Y(FE_RN_81_0),
	.A(FE_RN_58_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_107_0 (
	.Y(FE_RN_80_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_106_0 (
	.Y(FE_RN_79_0),
	.A(FE_RN_56_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M FE_RC_105_0 (
	.Y(FE_RN_78_0),
	.C(FE_RN_81_0),
	.B(FE_RN_80_0),
	.A(FE_RN_79_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_104_0 (
	.Y(FE_RN_77_0),
	.B(FE_RN_82_0),
	.A(FE_RN_78_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M FE_RC_103_0 (
	.Y(FE_RN_76_0),
	.A(FE_RN_77_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_102_0 (
	.Y(FE_RN_75_0),
	.C(FE_RN_84_0),
	.B(\u_div/SumTmp[5][0] ),
	.A(FE_RN_76_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B11X4M FE_RC_100_0 (
	.Y(\u_div/CryTmp[5][2] ),
	.C0(FE_RN_35_0),
	.B0(FE_RN_36_0),
	.A1N(FE_RN_42_0),
	.A0(FE_RN_30_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_99_0 (
	.Y(FE_RN_74_0),
	.A(FE_RN_42_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X3M FE_RC_98_0 (
	.Y(FE_RN_73_0),
	.B0(FE_RN_35_0),
	.A1(FE_RN_74_0),
	.A0(FE_RN_30_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_97_0 (
	.Y(FE_RN_72_0),
	.A(FE_RN_36_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_94_0 (
	.Y(FE_RN_69_0),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_92_0 (
	.Y(quotient[6]),
	.B(FE_RN_28_0),
	.A(FE_RN_31_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_91_0 (
	.Y(FE_RN_68_0),
	.A(FE_RN_56_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_90_0 (
	.Y(FE_RN_67_0),
	.A(FE_RN_58_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_89_0 (
	.Y(\u_div/PartRem[6][2] ),
	.B(FE_RN_68_0),
	.A(FE_RN_67_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_88_0 (
	.Y(FE_RN_66_0),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_87_0 (
	.Y(FE_RN_65_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M FE_RC_86_0 (
	.Y(FE_RN_64_0),
	.B1(\u_div/PartRem[7][1] ),
	.B0(FE_RN_65_0),
	.A1(n16),
	.A0(FE_RN_66_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_85_0 (
	.Y(FE_RN_63_0),
	.B(n16),
	.A(\u_div/SumTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X4M FE_RC_84_0 (
	.Y(FE_RN_62_0),
	.S0(FE_RN_57_0),
	.B(FE_RN_63_0),
	.A(FE_RN_64_0), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR2X2M FE_RC_83_0 (
	.Y(\u_div/SumTmp[5][2] ),
	.B(\u_div/CryTmp[5][2] ),
	.A(FE_RN_62_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_80_0 (
	.Y(FE_RN_59_0),
	.A(\u_div/PartRem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X8M FE_RC_79_0 (
	.Y(FE_RN_58_0),
	.B(FE_RN_59_0),
	.A(FE_RN_57_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X5M FE_RC_78_0 (
	.Y(FE_RN_57_0),
	.B(FE_RN_31_0),
	.A(FE_RN_28_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X8M FE_RC_77_0 (
	.Y(FE_RN_56_0),
	.B(\u_div/SumTmp[6][1] ),
	.A(FE_RN_57_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X6M FE_RC_76_0 (
	.Y(FE_RN_55_0),
	.B0(n16),
	.A1(FE_RN_56_0),
	.A0(FE_RN_58_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_74_0 (
	.Y(\u_div/PartRem[6][1] ),
	.S0(FE_RN_30_0),
	.B(FE_RN_33_0),
	.A(FE_RN_34_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_73_0 (
	.Y(FE_RN_54_0),
	.A(\u_div/CryTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_72_0 (
	.Y(FE_RN_53_0),
	.A(\u_div/CryTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_71_0 (
	.Y(FE_RN_52_0),
	.B(n17),
	.A(FE_RN_34_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X6M FE_RC_70_0 (
	.Y(FE_RN_51_0),
	.B0(FE_RN_52_0),
	.A1(n17),
	.A0(FE_RN_34_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X3M FE_RC_69_0 (
	.Y(FE_RN_50_0),
	.B(FE_RN_53_0),
	.A(FE_RN_51_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X4M FE_RC_68_0 (
	.Y(FE_RN_49_0),
	.B0(FE_RN_50_0),
	.A1(FE_RN_54_0),
	.A0(FE_RN_51_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_67_0 (
	.Y(FE_RN_48_0),
	.A(\u_div/CryTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_66_0 (
	.Y(FE_RN_47_0),
	.A(\u_div/CryTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M FE_RC_65_0 (
	.Y(FE_RN_46_0),
	.B(n17),
	.A(FE_RN_33_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB2X4M FE_RC_64_0 (
	.Y(FE_RN_45_0),
	.B1(FE_RN_46_0),
	.B0(FE_RN_47_0),
	.A1N(FE_RN_48_0),
	.A0N(FE_RN_46_0), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X2M FE_RC_63_0 (
	.Y(\u_div/SumTmp[5][1] ),
	.S0(FE_RN_30_0),
	.B(FE_RN_45_0),
	.A(FE_RN_49_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_62_0 (
	.Y(FE_RN_44_0),
	.A(FE_RN_34_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_61_0 (
	.Y(FE_RN_43_0),
	.A(FE_RN_39_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M FE_RC_60_0 (
	.Y(FE_RN_42_0),
	.B(FE_RN_43_0),
	.AN(FE_RN_44_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_59_0 (
	.Y(FE_RN_41_0),
	.A(\u_div/CryTmp[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_58_0 (
	.Y(FE_RN_40_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_57_0 (
	.Y(FE_RN_39_0),
	.B(FE_RN_41_0),
	.A(FE_RN_40_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_56_0 (
	.Y(FE_RN_38_0),
	.A(FE_RN_39_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M FE_RC_55_0 (
	.Y(FE_RN_37_0),
	.B(FE_RN_33_0),
	.A(FE_RN_38_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X3M FE_RC_54_0 (
	.Y(FE_RN_36_0),
	.B(FE_RN_30_0),
	.A(FE_RN_37_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M FE_RC_53_0 (
	.Y(FE_RN_35_0),
	.B(\u_div/CryTmp[5][1] ),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_50_0 (
	.Y(FE_RN_34_0),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_49_0 (
	.Y(FE_RN_33_0),
	.A(\u_div/SumTmp[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_48_0 (
	.Y(FE_RN_32_0),
	.A(FE_RN_14_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_47_0 (
	.Y(FE_RN_31_0),
	.C(FE_RN_27_0),
	.B(FE_RN_13_0),
	.AN(FE_RN_32_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_46_0 (
	.Y(FE_RN_30_0),
	.B(FE_RN_28_0),
	.A(FE_RN_31_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_44_0 (
	.Y(FE_RN_29_0),
	.A(FE_RN_17_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X3M FE_RC_43_0 (
	.Y(FE_RN_28_0),
	.C(FE_RN_29_0),
	.B(n16),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_42_0 (
	.Y(FE_RN_27_0),
	.B(n16),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_39_0 (
	.Y(\u_div/PartRem[7][1] ),
	.C(FE_RN_5_0),
	.B(FE_RN_9_0),
	.A(FE_RN_10_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_38_0 (
	.Y(FE_RN_25_0),
	.A(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_37_0 (
	.Y(FE_RN_24_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_36_0 (
	.Y(FE_RN_23_0),
	.A(FE_RN_18_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M FE_RC_35_0 (
	.Y(FE_RN_22_0),
	.B0(FE_RN_23_0),
	.A1N(FE_RN_24_0),
	.A0N(FE_RN_25_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_34_0 (
	.Y(FE_RN_21_0),
	.A(FE_RN_18_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M FE_RC_33_0 (
	.Y(FE_RN_20_0),
	.B(FE_RN_14_0),
	.A(FE_RN_21_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_32_0 (
	.Y(FE_RN_19_0),
	.B(FE_RN_13_0),
	.A(FE_RN_20_0), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X4M FE_RC_31_0 (
	.Y(\u_div/SumTmp[6][1] ),
	.B0(FE_RN_19_0),
	.A1(FE_RN_22_0),
	.A0(FE_RN_13_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_30_0 (
	.Y(FE_RN_18_0),
	.B(\u_div/CryTmp[6][1] ),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_29_0 (
	.Y(FE_RN_17_0),
	.A(FE_RN_18_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_28_0 (
	.Y(FE_RN_16_0),
	.A(\u_div/CryTmp[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_27_0 (
	.Y(FE_RN_15_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X4M FE_RC_26_0 (
	.Y(FE_RN_14_0),
	.B(FE_RN_16_0),
	.A(FE_RN_15_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X6M FE_RC_25_0 (
	.Y(FE_RN_13_0),
	.C(FE_RN_9_0),
	.B(FE_RN_10_0),
	.A(FE_RN_5_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_22_0 (
	.Y(FE_RN_11_0),
	.A(FE_RN_7_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_21_0 (
	.Y(quotient[7]),
	.B(n20),
	.A(FE_RN_11_0), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X4M FE_RC_20_0 (
	.Y(FE_RN_10_0),
	.B(a[7]),
	.A(FE_RN_7_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX8M FE_RC_19_0 (
	.Y(FE_RN_9_0),
	.B(a[7]),
	.AN(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X4M FE_RC_18_0 (
	.Y(FE_RN_8_0),
	.B(FE_RN_4_0),
	.A(FE_RN_2_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3BX4M FE_RC_17_0 (
	.Y(FE_RN_7_0),
	.C(\u_div/CryTmp[7][1] ),
	.B(FE_RN_8_0),
	.AN(FE_RN_3_0), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_16_0 (
	.Y(FE_RN_6_0),
	.A(FE_RN_7_0), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X4M FE_RC_15_0 (
	.Y(FE_RN_5_0),
	.C(n20),
	.B(\u_div/SumTmp[7][0] ),
	.A(FE_RN_6_0), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X6M FE_RC_13_0 (
	.Y(n20),
	.C(n13),
	.B(n14),
	.A(n21), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X4M FE_RC_12_0 (
	.Y(n19),
	.B(n15),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_11_0 (
	.Y(FE_RN_4_0),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_10_0 (
	.Y(FE_RN_3_0),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M FE_RC_9_0 (
	.Y(FE_RN_2_0),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX10M FE_RC_1_0 (
	.Y(n13),
	.A(b[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_5  (
	.CO(\u_div/CryTmp[0][6] ),
	.CI(\u_div/CryTmp[0][5] ),
	.B(n13),
	.A(\u_div/PartRem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_6  (
	.CO(\u_div/CryTmp[0][7] ),
	.CI(\u_div/CryTmp[0][6] ),
	.B(n140),
	.A(\u_div/PartRem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_7  (
	.CO(quotient[0]),
	.CI(\u_div/CryTmp[0][7] ),
	.B(n148),
	.A(\u_div/PartRem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_1  (
	.CO(\u_div/CryTmp[0][2] ),
	.CI(\u_div/CryTmp[0][1] ),
	.B(n17),
	.A(\u_div/PartRem[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_2  (
	.CO(\u_div/CryTmp[0][3] ),
	.CI(\u_div/CryTmp[0][2] ),
	.B(n16),
	.A(\u_div/PartRem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_3  (
	.CO(\u_div/CryTmp[0][4] ),
	.CI(\u_div/CryTmp[0][3] ),
	.B(n15),
	.A(\u_div/PartRem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX2M \u_div/u_fa_PartRem_0_0_4  (
	.CO(\u_div/CryTmp[0][5] ),
	.CI(\u_div/CryTmp[0][4] ),
	.B(n14),
	.A(\u_div/PartRem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFHX1M \u_div/u_fa_PartRem_0_1_6  (
	.S(\u_div/SumTmp[1][6] ),
	.CO(\u_div/CryTmp[1][7] ),
	.CI(\u_div/CryTmp[1][6] ),
	.B(n140),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX14M U1 (
	.Y(n18),
	.A(b[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U2 (
	.Y(\u_div/SumTmp[7][0] ),
	.B(a[7]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U3 (
	.Y(\u_div/SumTmp[6][0] ),
	.B(a[6]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(\u_div/SumTmp[5][0] ),
	.B(a[5]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(\u_div/SumTmp[4][0] ),
	.B(a[4]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(\u_div/SumTmp[3][0] ),
	.B(a[3]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(\u_div/SumTmp[2][0] ),
	.B(a[2]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X2M U8 (
	.Y(\u_div/CryTmp[7][1] ),
	.B(a[7]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(\u_div/SumTmp[1][0] ),
	.B(a[1]),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U10 (
	.Y(\u_div/CryTmp[5][1] ),
	.B(n3),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U11 (
	.Y(n3),
	.A(a[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U12 (
	.Y(n2),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U13 (
	.Y(\u_div/CryTmp[4][1] ),
	.B(n5),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U14 (
	.Y(n5),
	.A(a[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n4),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U16 (
	.Y(\u_div/CryTmp[3][1] ),
	.B(n7),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U17 (
	.Y(n7),
	.A(a[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n6),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U19 (
	.Y(\u_div/CryTmp[2][1] ),
	.B(n8),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n8),
	.A(a[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U21 (
	.Y(\u_div/CryTmp[1][1] ),
	.B(n9),
	.A(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n9),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U23 (
	.Y(\u_div/CryTmp[0][1] ),
	.B(n10),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n10),
	.A(a[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U25 (
	.Y(\u_div/CryTmp[6][1] ),
	.B(n1),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX2M U26 (
	.Y(n1),
	.A(a[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX14M U28 (
	.Y(n17),
	.A(b[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX12M U29 (
	.Y(n16),
	.A(b[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX12M U30 (
	.Y(n15),
	.A(b[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX14M U31 (
	.Y(n14),
	.A(b[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U34 (
	.Y(\u_div/PartRem[1][7] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][6] ),
	.A(\u_div/PartRem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U35 (
	.Y(\u_div/PartRem[2][6] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][5] ),
	.A(\u_div/PartRem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U36 (
	.Y(\u_div/PartRem[3][5] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][4] ),
	.A(\u_div/PartRem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U37 (
	.Y(\u_div/PartRem[4][4] ),
	.S0(quotient[4]),
	.B(\u_div/SumTmp[4][3] ),
	.A(\u_div/PartRem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X1M U38 (
	.Y(\u_div/PartRem[5][3] ),
	.S0(quotient[5]),
	.B(\u_div/SumTmp[5][2] ),
	.A(\u_div/PartRem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U41 (
	.Y(\u_div/PartRem[1][6] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][5] ),
	.A(\u_div/PartRem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U42 (
	.Y(\u_div/PartRem[2][5] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][4] ),
	.A(\u_div/PartRem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U43 (
	.Y(\u_div/PartRem[3][4] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][3] ),
	.A(\u_div/PartRem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U47 (
	.Y(\u_div/PartRem[1][5] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][4] ),
	.A(\u_div/PartRem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U48 (
	.Y(\u_div/PartRem[2][4] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][3] ),
	.A(\u_div/PartRem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U49 (
	.Y(\u_div/PartRem[3][3] ),
	.S0(quotient[3]),
	.B(\u_div/SumTmp[3][2] ),
	.A(\u_div/PartRem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U52 (
	.Y(\u_div/PartRem[1][4] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][3] ),
	.A(\u_div/PartRem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U53 (
	.Y(\u_div/PartRem[2][3] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][2] ),
	.A(\u_div/PartRem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U56 (
	.Y(\u_div/PartRem[1][3] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][2] ),
	.A(\u_div/PartRem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U57 (
	.Y(\u_div/PartRem[2][2] ),
	.S0(quotient[2]),
	.B(\u_div/SumTmp[2][1] ),
	.A(\u_div/PartRem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U59 (
	.Y(\u_div/PartRem[1][2] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][1] ),
	.A(\u_div/PartRem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX2X2M U61 (
	.Y(\u_div/PartRem[1][1] ),
	.S0(quotient[1]),
	.B(\u_div/SumTmp[1][0] ),
	.A(a[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X8M U70 (
	.Y(n21),
	.B(b[7]),
	.A(b[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X8M U71 (
	.Y(quotient[1]),
	.B(n148),
	.A(\u_div/CryTmp[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_sub_0 (
	A, 
	B, 
	CI, 
	DIFF, 
	CO, 
	n135, 
	n137, 
	n139, 
	n148, 
	n150, 
	n149, 
	n158, 
	n140, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] DIFF;
   output CO;
   input n135;
   input n137;
   input n139;
   input n148;
   input n150;
   input n149;
   input n158;
   input n140;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire [9:0] carry;

   // Module instantiations
   ADDFX2M U2_1 (
	.S(DIFF[1]),
	.CO(carry[2]),
	.CI(carry[1]),
	.B(n9),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_5 (
	.S(DIFF[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(n149),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_4 (
	.S(DIFF[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(n6),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_3 (
	.S(DIFF[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(n7),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_2 (
	.S(DIFF[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(n8),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_7 (
	.S(DIFF[7]),
	.CO(carry[8]),
	.CI(carry[7]),
	.B(n148),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U2_6 (
	.S(DIFF[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(n140),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U1 (
	.Y(DIFF[0]),
	.B(A[0]),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U2 (
	.Y(DIFF[8]),
	.A(carry[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U6 (
	.Y(n8),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U7 (
	.Y(n7),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n6),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U10 (
	.Y(carry[1]),
	.B(n1),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U11 (
	.Y(n9),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n1),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_add_0 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [8:0] A;
   input [8:0] B;
   input CI;
   output [8:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire [8:1] carry;

   // Module instantiations
   ADDFX2M U1_7 (
	.S(SUM[7]),
	.CO(SUM[8]),
	.CI(carry[7]),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_1 (
	.S(SUM[1]),
	.CO(carry[2]),
	.CI(n1),
	.B(B[1]),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_5 (
	.S(SUM[5]),
	.CO(carry[6]),
	.CI(carry[5]),
	.B(B[5]),
	.A(A[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_4 (
	.S(SUM[4]),
	.CO(carry[5]),
	.CI(carry[4]),
	.B(B[4]),
	.A(A[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_3 (
	.S(SUM[3]),
	.CO(carry[4]),
	.CI(carry[3]),
	.B(B[3]),
	.A(A[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_2 (
	.S(SUM[2]),
	.CO(carry[3]),
	.CI(carry[2]),
	.B(B[2]),
	.A(A[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M U1_6 (
	.S(SUM[6]),
	.CO(carry[7]),
	.CI(carry[6]),
	.B(B[6]),
	.A(A[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U1 (
	.Y(n1),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U2 (
	.Y(SUM[0]),
	.B(A[0]),
	.A(B[0]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW02_mult_0 (
	A, 
	B, 
	TC, 
	PRODUCT, 
	n135, 
	n137, 
	n139, 
	n158, 
	n157, 
	n156, 
	n155, 
	n154, 
	n153, 
	n152, 
	n151, 
	n148, 
	n149, 
	n140, 
	VDD, 
	VSS);
   input [7:0] A;
   input [7:0] B;
   input TC;
   output [15:0] PRODUCT;
   input n135;
   input n137;
   input n139;
   input n158;
   input n157;
   input n156;
   input n155;
   input n154;
   input n153;
   input n152;
   input n151;
   input n148;
   input n149;
   input n140;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \ab[7][7] ;
   wire \ab[7][6] ;
   wire \ab[7][5] ;
   wire \ab[7][4] ;
   wire \ab[7][3] ;
   wire \ab[7][2] ;
   wire \ab[7][1] ;
   wire \ab[7][0] ;
   wire \ab[6][7] ;
   wire \ab[6][6] ;
   wire \ab[6][5] ;
   wire \ab[6][4] ;
   wire \ab[6][3] ;
   wire \ab[6][2] ;
   wire \ab[6][1] ;
   wire \ab[6][0] ;
   wire \ab[5][7] ;
   wire \ab[5][6] ;
   wire \ab[5][5] ;
   wire \ab[5][4] ;
   wire \ab[5][3] ;
   wire \ab[5][2] ;
   wire \ab[5][1] ;
   wire \ab[5][0] ;
   wire \ab[4][7] ;
   wire \ab[4][6] ;
   wire \ab[4][5] ;
   wire \ab[4][4] ;
   wire \ab[4][3] ;
   wire \ab[4][2] ;
   wire \ab[4][1] ;
   wire \ab[4][0] ;
   wire \ab[3][7] ;
   wire \ab[3][6] ;
   wire \ab[3][5] ;
   wire \ab[3][4] ;
   wire \ab[3][3] ;
   wire \ab[3][2] ;
   wire \ab[3][1] ;
   wire \ab[3][0] ;
   wire \ab[2][7] ;
   wire \ab[2][6] ;
   wire \ab[2][5] ;
   wire \ab[2][4] ;
   wire \ab[2][3] ;
   wire \ab[2][2] ;
   wire \ab[2][1] ;
   wire \ab[2][0] ;
   wire \ab[1][7] ;
   wire \ab[1][6] ;
   wire \ab[1][5] ;
   wire \ab[1][4] ;
   wire \ab[1][3] ;
   wire \ab[1][2] ;
   wire \ab[1][1] ;
   wire \ab[1][0] ;
   wire \ab[0][7] ;
   wire \ab[0][6] ;
   wire \ab[0][5] ;
   wire \ab[0][4] ;
   wire \ab[0][3] ;
   wire \ab[0][2] ;
   wire \ab[0][1] ;
   wire \CARRYB[7][6] ;
   wire \CARRYB[7][5] ;
   wire \CARRYB[7][4] ;
   wire \CARRYB[7][3] ;
   wire \CARRYB[7][2] ;
   wire \CARRYB[7][1] ;
   wire \CARRYB[7][0] ;
   wire \CARRYB[6][6] ;
   wire \CARRYB[6][5] ;
   wire \CARRYB[6][4] ;
   wire \CARRYB[6][3] ;
   wire \CARRYB[6][2] ;
   wire \CARRYB[6][1] ;
   wire \CARRYB[6][0] ;
   wire \CARRYB[5][6] ;
   wire \CARRYB[5][5] ;
   wire \CARRYB[5][4] ;
   wire \CARRYB[5][3] ;
   wire \CARRYB[5][2] ;
   wire \CARRYB[5][1] ;
   wire \CARRYB[5][0] ;
   wire \CARRYB[4][6] ;
   wire \CARRYB[4][5] ;
   wire \CARRYB[4][4] ;
   wire \CARRYB[4][3] ;
   wire \CARRYB[4][2] ;
   wire \CARRYB[4][1] ;
   wire \CARRYB[4][0] ;
   wire \CARRYB[3][6] ;
   wire \CARRYB[3][5] ;
   wire \CARRYB[3][4] ;
   wire \CARRYB[3][3] ;
   wire \CARRYB[3][2] ;
   wire \CARRYB[3][1] ;
   wire \CARRYB[3][0] ;
   wire \CARRYB[2][6] ;
   wire \CARRYB[2][5] ;
   wire \CARRYB[2][4] ;
   wire \CARRYB[2][3] ;
   wire \CARRYB[2][2] ;
   wire \CARRYB[2][1] ;
   wire \CARRYB[2][0] ;
   wire \SUMB[7][6] ;
   wire \SUMB[7][5] ;
   wire \SUMB[7][4] ;
   wire \SUMB[7][3] ;
   wire \SUMB[7][2] ;
   wire \SUMB[7][1] ;
   wire \SUMB[7][0] ;
   wire \SUMB[6][6] ;
   wire \SUMB[6][5] ;
   wire \SUMB[6][4] ;
   wire \SUMB[6][3] ;
   wire \SUMB[6][2] ;
   wire \SUMB[6][1] ;
   wire \SUMB[5][6] ;
   wire \SUMB[5][5] ;
   wire \SUMB[5][4] ;
   wire \SUMB[5][3] ;
   wire \SUMB[5][2] ;
   wire \SUMB[5][1] ;
   wire \SUMB[4][6] ;
   wire \SUMB[4][5] ;
   wire \SUMB[4][4] ;
   wire \SUMB[4][3] ;
   wire \SUMB[4][2] ;
   wire \SUMB[4][1] ;
   wire \SUMB[3][6] ;
   wire \SUMB[3][5] ;
   wire \SUMB[3][4] ;
   wire \SUMB[3][3] ;
   wire \SUMB[3][2] ;
   wire \SUMB[3][1] ;
   wire \SUMB[2][6] ;
   wire \SUMB[2][5] ;
   wire \SUMB[2][4] ;
   wire \SUMB[2][3] ;
   wire \SUMB[2][2] ;
   wire \SUMB[2][1] ;
   wire \SUMB[1][6] ;
   wire \SUMB[1][5] ;
   wire \SUMB[1][4] ;
   wire \SUMB[1][3] ;
   wire \SUMB[1][2] ;
   wire \SUMB[1][1] ;
   wire \A1[12] ;
   wire \A1[11] ;
   wire \A1[10] ;
   wire \A1[9] ;
   wire \A1[8] ;
   wire \A1[7] ;
   wire \A1[6] ;
   wire \A1[4] ;
   wire \A1[3] ;
   wire \A1[2] ;
   wire \A1[1] ;
   wire \A1[0] ;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n38;
   wire n39;

   // Module instantiations
   ADDFX2M S1_6_0 (
	.S(\A1[4] ),
	.CO(\CARRYB[6][0] ),
	.CI(\SUMB[5][1] ),
	.B(\CARRYB[5][0] ),
	.A(\ab[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_5_0 (
	.S(\A1[3] ),
	.CO(\CARRYB[5][0] ),
	.CI(\SUMB[4][1] ),
	.B(\CARRYB[4][0] ),
	.A(\ab[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_4_0 (
	.S(\A1[2] ),
	.CO(\CARRYB[4][0] ),
	.CI(\SUMB[3][1] ),
	.B(\CARRYB[3][0] ),
	.A(\ab[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_3_0 (
	.S(\A1[1] ),
	.CO(\CARRYB[3][0] ),
	.CI(\SUMB[2][1] ),
	.B(\CARRYB[2][0] ),
	.A(\ab[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_5 (
	.S(\SUMB[6][5] ),
	.CO(\CARRYB[6][5] ),
	.CI(\SUMB[5][6] ),
	.B(\CARRYB[5][5] ),
	.A(\ab[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_4 (
	.S(\SUMB[6][4] ),
	.CO(\CARRYB[6][4] ),
	.CI(\SUMB[5][5] ),
	.B(\CARRYB[5][4] ),
	.A(\ab[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_5 (
	.S(\SUMB[5][5] ),
	.CO(\CARRYB[5][5] ),
	.CI(\SUMB[4][6] ),
	.B(\CARRYB[4][5] ),
	.A(\ab[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_3 (
	.S(\SUMB[6][3] ),
	.CO(\CARRYB[6][3] ),
	.CI(\SUMB[5][4] ),
	.B(\CARRYB[5][3] ),
	.A(\ab[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_4 (
	.S(\SUMB[5][4] ),
	.CO(\CARRYB[5][4] ),
	.CI(\SUMB[4][5] ),
	.B(\CARRYB[4][4] ),
	.A(\ab[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_1 (
	.S(\SUMB[6][1] ),
	.CO(\CARRYB[6][1] ),
	.CI(\SUMB[5][2] ),
	.B(\CARRYB[5][1] ),
	.A(\ab[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_6_2 (
	.S(\SUMB[6][2] ),
	.CO(\CARRYB[6][2] ),
	.CI(\SUMB[5][3] ),
	.B(\CARRYB[5][2] ),
	.A(\ab[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_5 (
	.S(\SUMB[4][5] ),
	.CO(\CARRYB[4][5] ),
	.CI(\SUMB[3][6] ),
	.B(\CARRYB[3][5] ),
	.A(\ab[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_1 (
	.S(\SUMB[5][1] ),
	.CO(\CARRYB[5][1] ),
	.CI(\SUMB[4][2] ),
	.B(\CARRYB[4][1] ),
	.A(\ab[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_2 (
	.S(\SUMB[5][2] ),
	.CO(\CARRYB[5][2] ),
	.CI(\SUMB[4][3] ),
	.B(\CARRYB[4][2] ),
	.A(\ab[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_5_3 (
	.S(\SUMB[5][3] ),
	.CO(\CARRYB[5][3] ),
	.CI(\SUMB[4][4] ),
	.B(\CARRYB[4][3] ),
	.A(\ab[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_1 (
	.S(\SUMB[4][1] ),
	.CO(\CARRYB[4][1] ),
	.CI(\SUMB[3][2] ),
	.B(\CARRYB[3][1] ),
	.A(\ab[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_2 (
	.S(\SUMB[4][2] ),
	.CO(\CARRYB[4][2] ),
	.CI(\SUMB[3][3] ),
	.B(\CARRYB[3][2] ),
	.A(\ab[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_3 (
	.S(\SUMB[4][3] ),
	.CO(\CARRYB[4][3] ),
	.CI(\SUMB[3][4] ),
	.B(\CARRYB[3][3] ),
	.A(\ab[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_4_4 (
	.S(\SUMB[4][4] ),
	.CO(\CARRYB[4][4] ),
	.CI(\SUMB[3][5] ),
	.B(\CARRYB[3][4] ),
	.A(\ab[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_1 (
	.S(\SUMB[3][1] ),
	.CO(\CARRYB[3][1] ),
	.CI(\SUMB[2][2] ),
	.B(\CARRYB[2][1] ),
	.A(\ab[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_2 (
	.S(\SUMB[3][2] ),
	.CO(\CARRYB[3][2] ),
	.CI(\SUMB[2][3] ),
	.B(\CARRYB[2][2] ),
	.A(\ab[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_3 (
	.S(\SUMB[3][3] ),
	.CO(\CARRYB[3][3] ),
	.CI(\SUMB[2][4] ),
	.B(\CARRYB[2][3] ),
	.A(\ab[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_4 (
	.S(\SUMB[3][4] ),
	.CO(\CARRYB[3][4] ),
	.CI(\SUMB[2][5] ),
	.B(\CARRYB[2][4] ),
	.A(\ab[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_3_5 (
	.S(\SUMB[3][5] ),
	.CO(\CARRYB[3][5] ),
	.CI(\SUMB[2][6] ),
	.B(\CARRYB[2][5] ),
	.A(\ab[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_6_6 (
	.S(\SUMB[6][6] ),
	.CO(\CARRYB[6][6] ),
	.CI(\ab[5][7] ),
	.B(\CARRYB[5][6] ),
	.A(\ab[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_5_6 (
	.S(\SUMB[5][6] ),
	.CO(\CARRYB[5][6] ),
	.CI(\ab[4][7] ),
	.B(\CARRYB[4][6] ),
	.A(\ab[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_4_6 (
	.S(\SUMB[4][6] ),
	.CO(\CARRYB[4][6] ),
	.CI(\ab[3][7] ),
	.B(\CARRYB[3][6] ),
	.A(\ab[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_3_6 (
	.S(\SUMB[3][6] ),
	.CO(\CARRYB[3][6] ),
	.CI(\ab[2][7] ),
	.B(\CARRYB[2][6] ),
	.A(\ab[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S3_2_6 (
	.S(\SUMB[2][6] ),
	.CO(\CARRYB[2][6] ),
	.CI(\ab[1][7] ),
	.B(n8),
	.A(\ab[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S1_2_0 (
	.S(\A1[0] ),
	.CO(\CARRYB[2][0] ),
	.CI(\SUMB[1][1] ),
	.B(n9),
	.A(\ab[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_1 (
	.S(\SUMB[2][1] ),
	.CO(\CARRYB[2][1] ),
	.CI(\SUMB[1][2] ),
	.B(n7),
	.A(\ab[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_2 (
	.S(\SUMB[2][2] ),
	.CO(\CARRYB[2][2] ),
	.CI(\SUMB[1][3] ),
	.B(n6),
	.A(\ab[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_3 (
	.S(\SUMB[2][3] ),
	.CO(\CARRYB[2][3] ),
	.CI(\SUMB[1][4] ),
	.B(n5),
	.A(\ab[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_4 (
	.S(\SUMB[2][4] ),
	.CO(\CARRYB[2][4] ),
	.CI(\SUMB[1][5] ),
	.B(n4),
	.A(\ab[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S2_2_5 (
	.S(\SUMB[2][5] ),
	.CO(\CARRYB[2][5] ),
	.CI(\SUMB[1][6] ),
	.B(n3),
	.A(\ab[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_0 (
	.S(\SUMB[7][0] ),
	.CO(\CARRYB[7][0] ),
	.CI(\SUMB[6][1] ),
	.B(\CARRYB[6][0] ),
	.A(\ab[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S5_6 (
	.S(\SUMB[7][6] ),
	.CO(\CARRYB[7][6] ),
	.CI(\ab[6][7] ),
	.B(\CARRYB[6][6] ),
	.A(\ab[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_5 (
	.S(\SUMB[7][5] ),
	.CO(\CARRYB[7][5] ),
	.CI(\SUMB[6][6] ),
	.B(\CARRYB[6][5] ),
	.A(\ab[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_4 (
	.S(\SUMB[7][4] ),
	.CO(\CARRYB[7][4] ),
	.CI(\SUMB[6][5] ),
	.B(\CARRYB[6][4] ),
	.A(\ab[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_3 (
	.S(\SUMB[7][3] ),
	.CO(\CARRYB[7][3] ),
	.CI(\SUMB[6][4] ),
	.B(\CARRYB[6][3] ),
	.A(\ab[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_2 (
	.S(\SUMB[7][2] ),
	.CO(\CARRYB[7][2] ),
	.CI(\SUMB[6][3] ),
	.B(\CARRYB[6][2] ),
	.A(\ab[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDFX2M S4_1 (
	.S(\SUMB[7][1] ),
	.CO(\CARRYB[7][1] ),
	.CI(\SUMB[6][2] ),
	.B(\CARRYB[6][1] ),
	.A(\ab[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U2 (
	.Y(n3),
	.B(\ab[1][5] ),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U3 (
	.Y(n4),
	.B(\ab[1][4] ),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(n5),
	.B(\ab[1][3] ),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U5 (
	.Y(n6),
	.B(\ab[1][2] ),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U6 (
	.Y(n7),
	.B(\ab[1][1] ),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U7 (
	.Y(n8),
	.B(\ab[1][6] ),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n9),
	.B(\ab[1][0] ),
	.A(\ab[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U9 (
	.Y(n10),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U10 (
	.Y(n22),
	.A(\ab[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U11 (
	.Y(\A1[7] ),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U12 (
	.Y(PRODUCT[1]),
	.B(\ab[0][1] ),
	.A(\ab[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(\A1[12] ),
	.B(\ab[7][7] ),
	.A(\CARRYB[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U14 (
	.Y(\A1[8] ),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U15 (
	.Y(\A1[10] ),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U16 (
	.Y(\A1[9] ),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U17 (
	.Y(\A1[11] ),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n23),
	.A(\ab[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n21),
	.A(\ab[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n20),
	.A(\ab[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U21 (
	.Y(n19),
	.A(\ab[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U22 (
	.Y(n18),
	.A(\ab[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U23 (
	.Y(n11),
	.B(\SUMB[7][1] ),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U24 (
	.Y(n17),
	.A(\SUMB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U25 (
	.Y(n12),
	.B(\SUMB[7][2] ),
	.A(\CARRYB[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U26 (
	.Y(n13),
	.B(\SUMB[7][4] ),
	.A(\CARRYB[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U27 (
	.Y(n14),
	.B(\SUMB[7][6] ),
	.A(\CARRYB[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U28 (
	.Y(n15),
	.B(\SUMB[7][3] ),
	.A(\CARRYB[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U29 (
	.Y(n16),
	.B(\SUMB[7][5] ),
	.A(\CARRYB[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U30 (
	.Y(\A1[6] ),
	.B(n17),
	.A(\CARRYB[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U31 (
	.Y(\SUMB[1][6] ),
	.B(n23),
	.A(\ab[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U32 (
	.Y(\SUMB[1][5] ),
	.B(n22),
	.A(\ab[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U33 (
	.Y(\SUMB[1][4] ),
	.B(n21),
	.A(\ab[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U34 (
	.Y(\SUMB[1][3] ),
	.B(n20),
	.A(\ab[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U35 (
	.Y(\SUMB[1][2] ),
	.B(n19),
	.A(\ab[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U36 (
	.Y(\SUMB[1][1] ),
	.B(n18),
	.A(\ab[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n38),
	.A(A[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n39),
	.A(A[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n29),
	.A(B[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U48 (
	.Y(n28),
	.A(B[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U50 (
	.Y(n27),
	.A(B[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U52 (
	.Y(n30),
	.A(B[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U54 (
	.Y(\ab[7][7] ),
	.B(n148),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U55 (
	.Y(\ab[7][6] ),
	.B(n140),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U56 (
	.Y(\ab[7][5] ),
	.B(n149),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U57 (
	.Y(\ab[7][4] ),
	.B(n27),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U58 (
	.Y(\ab[7][3] ),
	.B(n28),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U59 (
	.Y(\ab[7][2] ),
	.B(n29),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U60 (
	.Y(\ab[7][1] ),
	.B(n30),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U61 (
	.Y(\ab[7][0] ),
	.B(n135),
	.A(n151), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U62 (
	.Y(\ab[6][7] ),
	.B(n152),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U63 (
	.Y(\ab[6][6] ),
	.B(n152),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U64 (
	.Y(\ab[6][5] ),
	.B(n152),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U65 (
	.Y(\ab[6][4] ),
	.B(n152),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U66 (
	.Y(\ab[6][3] ),
	.B(n152),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U67 (
	.Y(\ab[6][2] ),
	.B(n152),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U68 (
	.Y(\ab[6][1] ),
	.B(n152),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U69 (
	.Y(\ab[6][0] ),
	.B(n152),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U70 (
	.Y(\ab[5][7] ),
	.B(n153),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U71 (
	.Y(\ab[5][6] ),
	.B(n153),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U72 (
	.Y(\ab[5][5] ),
	.B(n153),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U73 (
	.Y(\ab[5][4] ),
	.B(n153),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U74 (
	.Y(\ab[5][3] ),
	.B(n153),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U75 (
	.Y(\ab[5][2] ),
	.B(n153),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U76 (
	.Y(\ab[5][1] ),
	.B(n153),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U77 (
	.Y(\ab[5][0] ),
	.B(n153),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U78 (
	.Y(\ab[4][7] ),
	.B(n154),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U79 (
	.Y(\ab[4][6] ),
	.B(n154),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U80 (
	.Y(\ab[4][5] ),
	.B(n154),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U81 (
	.Y(\ab[4][4] ),
	.B(n154),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U82 (
	.Y(\ab[4][3] ),
	.B(n154),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U83 (
	.Y(\ab[4][2] ),
	.B(n154),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U84 (
	.Y(\ab[4][1] ),
	.B(n154),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U85 (
	.Y(\ab[4][0] ),
	.B(n154),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U86 (
	.Y(\ab[3][7] ),
	.B(n155),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U87 (
	.Y(\ab[3][6] ),
	.B(n155),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U88 (
	.Y(\ab[3][5] ),
	.B(n155),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U89 (
	.Y(\ab[3][4] ),
	.B(n155),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U90 (
	.Y(\ab[3][3] ),
	.B(n155),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U91 (
	.Y(\ab[3][2] ),
	.B(n155),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U92 (
	.Y(\ab[3][1] ),
	.B(n155),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U93 (
	.Y(\ab[3][0] ),
	.B(n155),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U94 (
	.Y(\ab[2][7] ),
	.B(n156),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U95 (
	.Y(\ab[2][6] ),
	.B(n156),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U96 (
	.Y(\ab[2][5] ),
	.B(n156),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U97 (
	.Y(\ab[2][4] ),
	.B(n156),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U98 (
	.Y(\ab[2][3] ),
	.B(n156),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U99 (
	.Y(\ab[2][2] ),
	.B(n156),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U100 (
	.Y(\ab[2][1] ),
	.B(n156),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U101 (
	.Y(\ab[2][0] ),
	.B(n156),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U102 (
	.Y(\ab[1][7] ),
	.B(n38),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U103 (
	.Y(\ab[1][6] ),
	.B(n38),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U104 (
	.Y(\ab[1][5] ),
	.B(n38),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U105 (
	.Y(\ab[1][4] ),
	.B(n38),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U106 (
	.Y(\ab[1][3] ),
	.B(n38),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U107 (
	.Y(\ab[1][2] ),
	.B(n38),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U108 (
	.Y(\ab[1][1] ),
	.B(n38),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U109 (
	.Y(\ab[1][0] ),
	.B(n38),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U110 (
	.Y(\ab[0][7] ),
	.B(n39),
	.A(n148), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U111 (
	.Y(\ab[0][6] ),
	.B(n39),
	.A(n140), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U112 (
	.Y(\ab[0][5] ),
	.B(n39),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U113 (
	.Y(\ab[0][4] ),
	.B(n39),
	.A(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U114 (
	.Y(\ab[0][3] ),
	.B(n39),
	.A(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U115 (
	.Y(\ab[0][2] ),
	.B(n39),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U116 (
	.Y(\ab[0][1] ),
	.B(n39),
	.A(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U117 (
	.Y(PRODUCT[0]),
	.B(n39),
	.A(n135), 
	.VDD(VDD), 
	.VSS(VSS));
   ALU_DW01_add_1 FS_1 (
	.A({ 1'b0,
		\A1[12] ,
		\A1[11] ,
		\A1[10] ,
		\A1[9] ,
		\A1[8] ,
		\A1[7] ,
		\A1[6] ,
		\SUMB[7][0] ,
		\A1[4] ,
		\A1[3] ,
		\A1[2] ,
		\A1[1] ,
		\A1[0]  }),
	.B({ n10,
		n14,
		n16,
		n13,
		n15,
		n12,
		n11,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0,
		1'b0 }),
	.CI(1'b0),
	.SUM({ PRODUCT[15],
		PRODUCT[14],
		PRODUCT[13],
		PRODUCT[12],
		PRODUCT[11],
		PRODUCT[10],
		PRODUCT[9],
		PRODUCT[8],
		PRODUCT[7],
		PRODUCT[6],
		PRODUCT[5],
		PRODUCT[4],
		PRODUCT[3],
		PRODUCT[2] }), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ALU_DW01_add_1 (
	A, 
	B, 
	CI, 
	SUM, 
	CO, 
	VDD, 
	VSS);
   input [13:0] A;
   input [13:0] B;
   input CI;
   output [13:0] SUM;
   output CO;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \A[5] ;
   wire \A[4] ;
   wire \A[3] ;
   wire \A[2] ;
   wire \A[1] ;
   wire \A[0] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;

   assign SUM[6] = A[6] ;
   assign SUM[5] = \A[5]  ;
   assign \A[5]  = A[5] ;
   assign SUM[4] = \A[4]  ;
   assign \A[4]  = A[4] ;
   assign SUM[3] = \A[3]  ;
   assign \A[3]  = A[3] ;
   assign SUM[2] = \A[2]  ;
   assign \A[2]  = A[2] ;
   assign SUM[1] = \A[1]  ;
   assign \A[1]  = A[1] ;
   assign SUM[0] = \A[0]  ;
   assign \A[0]  = A[0] ;

   // Module instantiations
   AOI21BX2M U2 (
	.Y(n1),
	.B0N(n12),
	.A1(A[12]),
	.A0(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U3 (
	.Y(n8),
	.B(B[7]),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U4 (
	.Y(SUM[7]),
	.B(n2),
	.A(A[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U5 (
	.Y(n2),
	.A(B[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U6 (
	.Y(SUM[13]),
	.B(n1),
	.A(B[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U7 (
	.Y(SUM[9]),
	.B(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U8 (
	.Y(n4),
	.B(n6),
	.A(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U9 (
	.Y(SUM[8]),
	.B(n8),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U10 (
	.Y(n7),
	.B(n10),
	.AN(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X1M U11 (
	.Y(n12),
	.B0(B[12]),
	.A1(n11),
	.A0(A[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U12 (
	.Y(SUM[12]),
	.C(n11),
	.B(A[12]),
	.A(B[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21BX1M U13 (
	.Y(n11),
	.B0N(n15),
	.A1(n14),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U14 (
	.Y(SUM[11]),
	.B(n16),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U15 (
	.Y(n16),
	.B(n13),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U16 (
	.Y(n13),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U17 (
	.Y(n15),
	.B(A[11]),
	.A(B[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U18 (
	.Y(n14),
	.B0(n19),
	.A1(n18),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U19 (
	.Y(SUM[10]),
	.B(n18),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2BB1X1M U20 (
	.Y(n18),
	.B0(n5),
	.A1N(n6),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U21 (
	.Y(n5),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U22 (
	.Y(n6),
	.B(A[9]),
	.A(B[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X1M U23 (
	.Y(n3),
	.B0(n10),
	.A1(n9),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U24 (
	.Y(n10),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U25 (
	.Y(n9),
	.B(A[8]),
	.A(B[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U26 (
	.Y(n20),
	.B(n19),
	.AN(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U27 (
	.Y(n19),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U28 (
	.Y(n17),
	.B(A[10]),
	.A(B[10]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module ASYNC_FIFO_DATA_WIDTH8_ADDR_WIDTH4_NUM_STAGES2_test_1 (
	wclk, 
	rclk, 
	wrst_n, 
	rrst_n, 
	W_INC, 
	R_INC, 
	wr_data, 
	FULL, 
	EMPTY, 
	rd_data, 
	test_si3, 
	test_si2, 
	test_si1, 
	test_so3, 
	test_so2, 
	test_so1, 
	test_se, 
	TX_CLK_M__L3_N1, 
	CLK_R_M__L5_N1, 
	CLK_R_M__L5_N2, 
	CLK_R_M__L5_N3, 
	CLK_R_M__L5_N4, 
	VDD, 
	VSS);
   input wclk;
   input rclk;
   input wrst_n;
   input rrst_n;
   input W_INC;
   input R_INC;
   input [7:0] wr_data;
   output FULL;
   output EMPTY;
   output [7:0] rd_data;
   input test_si3;
   input test_si2;
   input test_si1;
   output test_so3;
   output test_so2;
   output test_so1;
   input test_se;
   input TX_CLK_M__L3_N1;
   input CLK_R_M__L5_N1;
   input CLK_R_M__L5_N2;
   input CLK_R_M__L5_N3;
   input CLK_R_M__L5_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN2_RST_SYNC_1_mux;
   wire n1;
   wire [3:0] waddr;
   wire [3:0] raddr;
   wire [4:0] wptr_async;
   wire [4:0] rq2_wptr_sync;
   wire [4:0] rptr_async;
   wire [4:0] wq2_rptr_sync;

   assign test_so2 = raddr[0] ;
   assign test_so3 = wptr_async[4] ;

   // Module instantiations
   CLKBUFX8M FE_OFC2_RST_SYNC_1_mux (
	.Y(FE_OFN2_RST_SYNC_1_mux),
	.A(wrst_n), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_MEM_CNTRL_DATA_WIDTH8_ADDR_WIDTH4_test_1 fifo_mem_cntrl (
	.i_w_clk(wclk),
	.i_rst_n(wrst_n),
	.i_w_inc(W_INC),
	.i_w_full(FULL),
	.i_wr_data({ wr_data[7],
		wr_data[6],
		wr_data[5],
		wr_data[4],
		wr_data[3],
		wr_data[2],
		wr_data[1],
		wr_data[0] }),
	.i_wr_addr({ waddr[3],
		waddr[2],
		waddr[1],
		waddr[0] }),
	.i_rd_addr({ raddr[3],
		raddr[2],
		raddr[1],
		raddr[0] }),
	.o_rd_data({ rd_data[7],
		rd_data[6],
		rd_data[5],
		rd_data[4],
		rd_data[3],
		rd_data[2],
		rd_data[1],
		rd_data[0] }),
	.test_si2(test_si2),
	.test_si1(rq2_wptr_sync[4]),
	.test_so2(n1),
	.test_so1(test_so1),
	.test_se(test_se),
	.FE_OFN2_RST_SYNC_1_mux(FE_OFN2_RST_SYNC_1_mux),
	.CLK_R_M__L5_N1(CLK_R_M__L5_N1),
	.CLK_R_M__L5_N2(CLK_R_M__L5_N2),
	.CLK_R_M__L5_N3(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   DF_SYNC_ADDR_WIDTH4_test_1 bit_sync_waddr (
	.i_clk(rclk),
	.i_rst_n(rrst_n),
	.i_r_d_ptr({ wptr_async[4],
		wptr_async[3],
		wptr_async[2],
		wptr_async[1],
		wptr_async[0] }),
	.wq2_r_d_ptr({ rq2_wptr_sync[4],
		rq2_wptr_sync[3],
		rq2_wptr_sync[2],
		rq2_wptr_sync[1],
		rq2_wptr_sync[0] }),
	.test_si(wq2_rptr_sync[4]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DF_SYNC_ADDR_WIDTH4_test_0 bit_sync_raddr (
	.i_clk(CLK_R_M__L5_N3),
	.i_rst_n(wrst_n),
	.i_r_d_ptr({ rptr_async[4],
		rptr_async[3],
		rptr_async[2],
		rptr_async[1],
		rptr_async[0] }),
	.wq2_r_d_ptr({ wq2_rptr_sync[4],
		wq2_rptr_sync[3],
		wq2_rptr_sync[2],
		wq2_rptr_sync[1],
		wq2_rptr_sync[0] }),
	.test_si(test_si1),
	.test_se(test_se),
	.CLK_R_M__L5_N4(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_RD_DATA_WIDTH8_ADDR_WIDTH4_test_1 fifo_rd (
	.i_r_clk(rclk),
	.i_rst_n(rrst_n),
	.i_r_inc(R_INC),
	.rq2_wptr({ rq2_wptr_sync[4],
		rq2_wptr_sync[3],
		rq2_wptr_sync[2],
		rq2_wptr_sync[1],
		rq2_wptr_sync[0] }),
	.o_r_empty(EMPTY),
	.o_rd_addr({ raddr[3],
		raddr[2],
		raddr[1],
		raddr[0] }),
	.o_rptr({ rptr_async[4],
		rptr_async[3],
		rptr_async[2],
		rptr_async[1],
		rptr_async[0] }),
	.test_si2(test_si3),
	.test_si1(n1),
	.test_se(test_se),
	.TX_CLK_M__L3_N1(TX_CLK_M__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   FIFO_WR_DATA_WIDTH8_ADDR_WIDTH4_test_1 fifo_wr (
	.i_w_clk(CLK_R_M__L5_N1),
	.i_rst_n(wrst_n),
	.i_w_inc(W_INC),
	.wq2_rptr({ wq2_rptr_sync[4],
		wq2_rptr_sync[3],
		wq2_rptr_sync[2],
		wq2_rptr_sync[1],
		wq2_rptr_sync[0] }),
	.o_w_full(FULL),
	.o_wr_addr({ waddr[3],
		waddr[2],
		waddr[1],
		waddr[0] }),
	.o_wptr({ wptr_async[4],
		wptr_async[3],
		wptr_async[2],
		wptr_async[1],
		wptr_async[0] }),
	.test_si(rptr_async[4]),
	.test_se(test_se),
	.FE_OFN2_RST_SYNC_1_mux(FE_OFN2_RST_SYNC_1_mux),
	.CLK_R_M__L5_N3(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_MEM_CNTRL_DATA_WIDTH8_ADDR_WIDTH4_test_1 (
	i_w_clk, 
	i_rst_n, 
	i_w_inc, 
	i_w_full, 
	i_wr_data, 
	i_wr_addr, 
	i_rd_addr, 
	o_rd_data, 
	test_si2, 
	test_si1, 
	test_so2, 
	test_so1, 
	test_se, 
	FE_OFN2_RST_SYNC_1_mux, 
	CLK_R_M__L5_N1, 
	CLK_R_M__L5_N2, 
	CLK_R_M__L5_N3, 
	VDD, 
	VSS);
   input i_w_clk;
   input i_rst_n;
   input i_w_inc;
   input i_w_full;
   input [7:0] i_wr_data;
   input [3:0] i_wr_addr;
   input [3:0] i_rd_addr;
   output [7:0] o_rd_data;
   input test_si2;
   input test_si1;
   output test_so2;
   output test_so1;
   input test_se;
   input FE_OFN2_RST_SYNC_1_mux;
   input CLK_R_M__L5_N1;
   input CLK_R_M__L5_N2;
   input CLK_R_M__L5_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire FE_OFN3_RST_SYNC_1_mux;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire \mem[0][7] ;
   wire \mem[0][6] ;
   wire \mem[0][5] ;
   wire \mem[0][4] ;
   wire \mem[0][3] ;
   wire \mem[0][2] ;
   wire \mem[0][1] ;
   wire \mem[0][0] ;
   wire \mem[1][7] ;
   wire \mem[1][6] ;
   wire \mem[1][5] ;
   wire \mem[1][4] ;
   wire \mem[1][3] ;
   wire \mem[1][2] ;
   wire \mem[1][1] ;
   wire \mem[1][0] ;
   wire \mem[2][7] ;
   wire \mem[2][6] ;
   wire \mem[2][5] ;
   wire \mem[2][4] ;
   wire \mem[2][3] ;
   wire \mem[2][2] ;
   wire \mem[2][1] ;
   wire \mem[2][0] ;
   wire \mem[3][7] ;
   wire \mem[3][6] ;
   wire \mem[3][5] ;
   wire \mem[3][4] ;
   wire \mem[3][3] ;
   wire \mem[3][2] ;
   wire \mem[3][1] ;
   wire \mem[3][0] ;
   wire \mem[4][7] ;
   wire \mem[4][6] ;
   wire \mem[4][5] ;
   wire \mem[4][4] ;
   wire \mem[4][3] ;
   wire \mem[4][2] ;
   wire \mem[4][1] ;
   wire \mem[4][0] ;
   wire \mem[5][7] ;
   wire \mem[5][6] ;
   wire \mem[5][5] ;
   wire \mem[5][4] ;
   wire \mem[5][3] ;
   wire \mem[5][2] ;
   wire \mem[5][1] ;
   wire \mem[5][0] ;
   wire \mem[6][7] ;
   wire \mem[6][6] ;
   wire \mem[6][5] ;
   wire \mem[6][4] ;
   wire \mem[6][3] ;
   wire \mem[6][2] ;
   wire \mem[6][1] ;
   wire \mem[6][0] ;
   wire \mem[7][7] ;
   wire \mem[7][6] ;
   wire \mem[7][5] ;
   wire \mem[7][4] ;
   wire \mem[7][3] ;
   wire \mem[7][2] ;
   wire \mem[7][1] ;
   wire \mem[7][0] ;
   wire \mem[8][7] ;
   wire \mem[8][6] ;
   wire \mem[8][5] ;
   wire \mem[8][4] ;
   wire \mem[8][3] ;
   wire \mem[8][2] ;
   wire \mem[8][1] ;
   wire \mem[8][0] ;
   wire \mem[9][7] ;
   wire \mem[9][6] ;
   wire \mem[9][5] ;
   wire \mem[9][4] ;
   wire \mem[9][3] ;
   wire \mem[9][2] ;
   wire \mem[9][1] ;
   wire \mem[9][0] ;
   wire \mem[10][7] ;
   wire \mem[10][6] ;
   wire \mem[10][5] ;
   wire \mem[10][4] ;
   wire \mem[10][3] ;
   wire \mem[10][2] ;
   wire \mem[10][1] ;
   wire \mem[10][0] ;
   wire \mem[11][7] ;
   wire \mem[11][6] ;
   wire \mem[11][5] ;
   wire \mem[11][4] ;
   wire \mem[11][3] ;
   wire \mem[11][2] ;
   wire \mem[11][1] ;
   wire \mem[11][0] ;
   wire \mem[12][7] ;
   wire \mem[12][6] ;
   wire \mem[12][5] ;
   wire \mem[12][4] ;
   wire \mem[12][3] ;
   wire \mem[12][2] ;
   wire \mem[12][1] ;
   wire \mem[12][0] ;
   wire \mem[13][7] ;
   wire \mem[13][6] ;
   wire \mem[13][5] ;
   wire \mem[13][4] ;
   wire \mem[13][3] ;
   wire \mem[13][2] ;
   wire \mem[13][1] ;
   wire \mem[13][0] ;
   wire \mem[14][7] ;
   wire \mem[14][6] ;
   wire \mem[14][5] ;
   wire \mem[14][4] ;
   wire \mem[14][3] ;
   wire \mem[14][2] ;
   wire \mem[14][1] ;
   wire \mem[14][0] ;
   wire \mem[15][7] ;
   wire \mem[15][6] ;
   wire \mem[15][5] ;
   wire \mem[15][4] ;
   wire \mem[15][3] ;
   wire \mem[15][2] ;
   wire \mem[15][1] ;
   wire \mem[15][0] ;
   wire n140;
   wire n141;
   wire n142;
   wire n143;
   wire n144;
   wire n145;
   wire n146;
   wire n147;
   wire n148;
   wire n149;
   wire n150;
   wire n151;
   wire n152;
   wire n153;
   wire n154;
   wire n155;
   wire n156;
   wire n157;
   wire n158;
   wire n159;
   wire n160;
   wire n161;
   wire n162;
   wire n163;
   wire n164;
   wire n165;
   wire n166;
   wire n167;
   wire n168;
   wire n169;
   wire n170;
   wire n171;
   wire n172;
   wire n173;
   wire n174;
   wire n175;
   wire n176;
   wire n177;
   wire n178;
   wire n179;
   wire n180;
   wire n181;
   wire n182;
   wire n183;
   wire n184;
   wire n185;
   wire n186;
   wire n187;
   wire n188;
   wire n189;
   wire n190;
   wire n191;
   wire n192;
   wire n193;
   wire n194;
   wire n195;
   wire n196;
   wire n197;
   wire n198;
   wire n199;
   wire n200;
   wire n201;
   wire n202;
   wire n203;
   wire n204;
   wire n205;
   wire n206;
   wire n207;
   wire n208;
   wire n209;
   wire n210;
   wire n211;
   wire n212;
   wire n213;
   wire n214;
   wire n215;
   wire n216;
   wire n217;
   wire n218;
   wire n219;
   wire n220;
   wire n221;
   wire n222;
   wire n223;
   wire n224;
   wire n225;
   wire n226;
   wire n227;
   wire n228;
   wire n229;
   wire n230;
   wire n231;
   wire n232;
   wire n233;
   wire n234;
   wire n235;
   wire n236;
   wire n237;
   wire n238;
   wire n239;
   wire n240;
   wire n241;
   wire n242;
   wire n243;
   wire n244;
   wire n245;
   wire n246;
   wire n247;
   wire n248;
   wire n249;
   wire n250;
   wire n251;
   wire n252;
   wire n253;
   wire n254;
   wire n255;
   wire n256;
   wire n257;
   wire n258;
   wire n259;
   wire n260;
   wire n261;
   wire n262;
   wire n263;
   wire n264;
   wire n265;
   wire n266;
   wire n267;
   wire n268;
   wire n269;
   wire n270;
   wire n271;
   wire n272;
   wire n273;
   wire n274;
   wire n275;
   wire n276;
   wire n277;
   wire n278;
   wire n279;
   wire n280;
   wire n281;
   wire n282;
   wire n283;
   wire n284;
   wire n285;
   wire n286;
   wire n287;
   wire n288;
   wire n289;
   wire n290;
   wire n291;
   wire n292;
   wire n293;
   wire n294;
   wire n129;
   wire n130;
   wire n131;
   wire n132;
   wire n133;
   wire n134;
   wire n135;
   wire n136;
   wire n137;
   wire n138;
   wire n139;
   wire n295;
   wire n296;
   wire n297;
   wire n298;
   wire n299;
   wire n300;
   wire n301;
   wire n302;
   wire n303;
   wire n304;
   wire n305;
   wire n306;
   wire n307;
   wire n308;
   wire n309;
   wire n310;
   wire n311;
   wire n312;
   wire n313;
   wire n314;
   wire n315;
   wire n316;
   wire n318;
   wire n319;
   wire n321;
   wire n322;
   wire n340;
   wire n341;
   wire n342;
   wire n343;
   wire n344;
   wire n345;
   wire n346;
   wire n347;
   wire n348;
   wire n349;
   wire n350;
   wire n354;
   wire n355;
   wire n356;
   wire n357;

   assign N10 = i_rd_addr[0] ;
   assign N11 = i_rd_addr[1] ;
   assign N12 = i_rd_addr[2] ;
   assign N13 = i_rd_addr[3] ;
   assign test_so1 = \mem[5][5]  ;
   assign test_so2 = \mem[15][7]  ;

   // Module instantiations
   BUFX8M FE_OFC3_RST_SYNC_1_mux (
	.Y(FE_OFN3_RST_SYNC_1_mux),
	.A(FE_OFN2_RST_SYNC_1_mux), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][7]  (
	.SI(\mem[1][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[1][7] ),
	.D(n286),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][6]  (
	.SI(\mem[1][5] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[1][6] ),
	.D(n285),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][5]  (
	.SI(\mem[1][4] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[1][5] ),
	.D(n284),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][4]  (
	.SI(\mem[1][3] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[1][4] ),
	.D(n283),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][3]  (
	.SI(\mem[1][2] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[1][3] ),
	.D(n282),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][2]  (
	.SI(\mem[1][1] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[1][2] ),
	.D(n281),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][1]  (
	.SI(\mem[1][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[1][1] ),
	.D(n280),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[1][0]  (
	.SI(\mem[0][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[1][0] ),
	.D(n279),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][7]  (
	.SI(\mem[5][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[5][7] ),
	.D(n254),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][6]  (
	.SI(test_si2),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[5][6] ),
	.D(n253),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][5]  (
	.SI(\mem[5][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[5][5] ),
	.D(n252),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][4]  (
	.SI(\mem[5][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[5][4] ),
	.D(n251),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][3]  (
	.SI(\mem[5][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[5][3] ),
	.D(n250),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][2]  (
	.SI(\mem[5][1] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[5][2] ),
	.D(n249),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][1]  (
	.SI(\mem[5][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[5][1] ),
	.D(n248),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[5][0]  (
	.SI(\mem[4][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[5][0] ),
	.D(n247),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][7]  (
	.SI(\mem[9][6] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[9][7] ),
	.D(n222),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][6]  (
	.SI(\mem[9][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[9][6] ),
	.D(n221),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][5]  (
	.SI(\mem[9][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[9][5] ),
	.D(n220),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][4]  (
	.SI(\mem[9][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[9][4] ),
	.D(n219),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][3]  (
	.SI(\mem[9][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[9][3] ),
	.D(n218),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][2]  (
	.SI(\mem[9][1] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[9][2] ),
	.D(n217),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][1]  (
	.SI(\mem[9][0] ),
	.SE(n356),
	.RN(i_rst_n),
	.Q(\mem[9][1] ),
	.D(n216),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[9][0]  (
	.SI(\mem[8][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[9][0] ),
	.D(n215),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][7]  (
	.SI(\mem[13][6] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[13][7] ),
	.D(n190),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][6]  (
	.SI(\mem[13][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[13][6] ),
	.D(n189),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][5]  (
	.SI(\mem[13][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[13][5] ),
	.D(n188),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][4]  (
	.SI(\mem[13][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[13][4] ),
	.D(n187),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][3]  (
	.SI(\mem[13][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[13][3] ),
	.D(n186),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][2]  (
	.SI(\mem[13][1] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[13][2] ),
	.D(n185),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][1]  (
	.SI(\mem[13][0] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[13][1] ),
	.D(n184),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[13][0]  (
	.SI(\mem[12][7] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[13][0] ),
	.D(n183),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][7]  (
	.SI(\mem[3][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[3][7] ),
	.D(n270),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][6]  (
	.SI(\mem[3][5] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[3][6] ),
	.D(n269),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][5]  (
	.SI(\mem[3][4] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[3][5] ),
	.D(n268),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][4]  (
	.SI(\mem[3][3] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[3][4] ),
	.D(n267),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][3]  (
	.SI(\mem[3][2] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[3][3] ),
	.D(n266),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][2]  (
	.SI(\mem[3][1] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[3][2] ),
	.D(n265),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][1]  (
	.SI(\mem[3][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[3][1] ),
	.D(n264),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[3][0]  (
	.SI(\mem[2][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[3][0] ),
	.D(n263),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][7]  (
	.SI(\mem[7][6] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[7][7] ),
	.D(n238),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][6]  (
	.SI(\mem[7][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[7][6] ),
	.D(n237),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][5]  (
	.SI(\mem[7][4] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[7][5] ),
	.D(n236),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][4]  (
	.SI(\mem[7][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[7][4] ),
	.D(n235),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][3]  (
	.SI(\mem[7][2] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[7][3] ),
	.D(n234),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][2]  (
	.SI(\mem[7][1] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[7][2] ),
	.D(n233),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][1]  (
	.SI(\mem[7][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[7][1] ),
	.D(n232),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[7][0]  (
	.SI(\mem[6][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[7][0] ),
	.D(n231),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][7]  (
	.SI(\mem[11][6] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[11][7] ),
	.D(n206),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][6]  (
	.SI(\mem[11][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[11][6] ),
	.D(n205),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][5]  (
	.SI(\mem[11][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[11][5] ),
	.D(n204),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][4]  (
	.SI(\mem[11][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[11][4] ),
	.D(n203),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][3]  (
	.SI(\mem[11][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[11][3] ),
	.D(n202),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][2]  (
	.SI(\mem[11][1] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[11][2] ),
	.D(n201),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][1]  (
	.SI(\mem[11][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[11][1] ),
	.D(n200),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[11][0]  (
	.SI(\mem[10][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[11][0] ),
	.D(n199),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][7]  (
	.SI(\mem[15][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[15][7] ),
	.D(n174),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][6]  (
	.SI(\mem[15][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[15][6] ),
	.D(n173),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][5]  (
	.SI(\mem[15][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[15][5] ),
	.D(n172),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][4]  (
	.SI(\mem[15][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[15][4] ),
	.D(n171),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][3]  (
	.SI(\mem[15][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[15][3] ),
	.D(n170),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][2]  (
	.SI(\mem[15][1] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[15][2] ),
	.D(n169),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][1]  (
	.SI(\mem[15][0] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[15][1] ),
	.D(n168),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[15][0]  (
	.SI(\mem[14][7] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[15][0] ),
	.D(n167),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][7]  (
	.SI(\mem[2][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[2][7] ),
	.D(n278),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][6]  (
	.SI(\mem[2][5] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[2][6] ),
	.D(n277),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][5]  (
	.SI(\mem[2][4] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[2][5] ),
	.D(n276),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][4]  (
	.SI(\mem[2][3] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[2][4] ),
	.D(n275),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][3]  (
	.SI(\mem[2][2] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[2][3] ),
	.D(n274),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][2]  (
	.SI(\mem[2][1] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[2][2] ),
	.D(n273),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][1]  (
	.SI(\mem[2][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[2][1] ),
	.D(n272),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[2][0]  (
	.SI(\mem[1][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[2][0] ),
	.D(n271),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][7]  (
	.SI(\mem[6][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[6][7] ),
	.D(n246),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][6]  (
	.SI(\mem[6][5] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[6][6] ),
	.D(n245),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][5]  (
	.SI(\mem[6][4] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[6][5] ),
	.D(n244),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][4]  (
	.SI(\mem[6][3] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[6][4] ),
	.D(n243),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][3]  (
	.SI(\mem[6][2] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[6][3] ),
	.D(n242),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][2]  (
	.SI(\mem[6][1] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[6][2] ),
	.D(n241),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][1]  (
	.SI(\mem[6][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[6][1] ),
	.D(n240),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[6][0]  (
	.SI(\mem[5][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[6][0] ),
	.D(n239),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][7]  (
	.SI(\mem[10][6] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[10][7] ),
	.D(n214),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][6]  (
	.SI(\mem[10][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[10][6] ),
	.D(n213),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][5]  (
	.SI(\mem[10][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[10][5] ),
	.D(n212),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][4]  (
	.SI(\mem[10][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[10][4] ),
	.D(n211),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][3]  (
	.SI(\mem[10][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[10][3] ),
	.D(n210),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][2]  (
	.SI(\mem[10][1] ),
	.SE(n357),
	.RN(i_rst_n),
	.Q(\mem[10][2] ),
	.D(n209),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][1]  (
	.SI(\mem[10][0] ),
	.SE(n356),
	.RN(i_rst_n),
	.Q(\mem[10][1] ),
	.D(n208),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[10][0]  (
	.SI(\mem[9][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[10][0] ),
	.D(n207),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][7]  (
	.SI(\mem[14][6] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[14][7] ),
	.D(n182),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][6]  (
	.SI(\mem[14][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[14][6] ),
	.D(n181),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][5]  (
	.SI(\mem[14][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[14][5] ),
	.D(n180),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][4]  (
	.SI(\mem[14][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[14][4] ),
	.D(n179),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][3]  (
	.SI(\mem[14][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[14][3] ),
	.D(n178),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][2]  (
	.SI(\mem[14][1] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[14][2] ),
	.D(n177),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][1]  (
	.SI(\mem[14][0] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[14][1] ),
	.D(n176),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[14][0]  (
	.SI(\mem[13][7] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[14][0] ),
	.D(n175),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][7]  (
	.SI(\mem[0][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[0][7] ),
	.D(n294),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][6]  (
	.SI(\mem[0][5] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[0][6] ),
	.D(n293),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][5]  (
	.SI(\mem[0][4] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[0][5] ),
	.D(n292),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][4]  (
	.SI(\mem[0][3] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[0][4] ),
	.D(n291),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][3]  (
	.SI(\mem[0][2] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[0][3] ),
	.D(n290),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][2]  (
	.SI(\mem[0][1] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[0][2] ),
	.D(n289),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][1]  (
	.SI(\mem[0][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[0][1] ),
	.D(n288),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[0][0]  (
	.SI(test_si1),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[0][0] ),
	.D(n287),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][7]  (
	.SI(\mem[4][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[4][7] ),
	.D(n262),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][6]  (
	.SI(\mem[4][5] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[4][6] ),
	.D(n261),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][5]  (
	.SI(\mem[4][4] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[4][5] ),
	.D(n260),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][4]  (
	.SI(\mem[4][3] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[4][4] ),
	.D(n259),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][3]  (
	.SI(\mem[4][2] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[4][3] ),
	.D(n258),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][2]  (
	.SI(\mem[4][1] ),
	.SE(n357),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[4][2] ),
	.D(n257),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][1]  (
	.SI(\mem[4][0] ),
	.SE(n356),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[4][1] ),
	.D(n256),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[4][0]  (
	.SI(\mem[3][7] ),
	.SE(n355),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[4][0] ),
	.D(n255),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][7]  (
	.SI(\mem[8][6] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[8][7] ),
	.D(n230),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][6]  (
	.SI(\mem[8][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[8][6] ),
	.D(n229),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][5]  (
	.SI(\mem[8][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[8][5] ),
	.D(n228),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][4]  (
	.SI(\mem[8][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[8][4] ),
	.D(n227),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][3]  (
	.SI(\mem[8][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[8][3] ),
	.D(n226),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][2]  (
	.SI(\mem[8][1] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[8][2] ),
	.D(n225),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][1]  (
	.SI(\mem[8][0] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[8][1] ),
	.D(n224),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[8][0]  (
	.SI(\mem[7][7] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[8][0] ),
	.D(n223),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][7]  (
	.SI(\mem[12][6] ),
	.SE(n354),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(\mem[12][7] ),
	.D(n198),
	.CK(CLK_R_M__L5_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][6]  (
	.SI(\mem[12][5] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[12][6] ),
	.D(n197),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][5]  (
	.SI(\mem[12][4] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[12][5] ),
	.D(n196),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][4]  (
	.SI(\mem[12][3] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[12][4] ),
	.D(n195),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][3]  (
	.SI(\mem[12][2] ),
	.SE(n354),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[12][3] ),
	.D(n194),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][2]  (
	.SI(\mem[12][1] ),
	.SE(n357),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[12][2] ),
	.D(n193),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][1]  (
	.SI(\mem[12][0] ),
	.SE(n356),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[12][1] ),
	.D(n192),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \mem_reg[12][0]  (
	.SI(\mem[11][7] ),
	.SE(n355),
	.RN(FE_OFN3_RST_SYNC_1_mux),
	.Q(\mem[12][0] ),
	.D(n191),
	.CK(CLK_R_M__L5_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U130 (
	.Y(n141),
	.B(n349),
	.A(n350), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U131 (
	.Y(n340),
	.A(i_wr_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U132 (
	.Y(n341),
	.A(i_wr_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U133 (
	.Y(n342),
	.A(i_wr_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U134 (
	.Y(n343),
	.A(i_wr_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U135 (
	.Y(n344),
	.A(i_wr_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U136 (
	.Y(n345),
	.A(i_wr_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U137 (
	.Y(n346),
	.A(i_wr_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U138 (
	.Y(n347),
	.A(i_wr_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U139 (
	.Y(n149),
	.B(i_wr_addr[2]),
	.A(n349), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U140 (
	.Y(n152),
	.B(i_wr_addr[2]),
	.A(i_wr_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U141 (
	.Y(n146),
	.B(i_wr_addr[1]),
	.A(n350), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U142 (
	.Y(n321),
	.A(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX4M U154 (
	.Y(n322),
	.A(n319), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U160 (
	.Y(n143),
	.B(n141),
	.A(n144), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U161 (
	.Y(n158),
	.B(n141),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX3M U162 (
	.Y(n318),
	.A(n316), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U163 (
	.Y(n319),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U166 (
	.Y(n145),
	.B(n142),
	.A(n146), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U167 (
	.Y(n147),
	.B(n144),
	.A(n146), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U168 (
	.Y(n148),
	.B(n142),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U169 (
	.Y(n150),
	.B(n144),
	.A(n149), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U170 (
	.Y(n151),
	.B(n142),
	.A(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U171 (
	.Y(n154),
	.B(n144),
	.A(n152), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U172 (
	.Y(n160),
	.B(n146),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U173 (
	.Y(n161),
	.B(n146),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U174 (
	.Y(n162),
	.B(n149),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U175 (
	.Y(n163),
	.B(n149),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U176 (
	.Y(n164),
	.B(n152),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U177 (
	.Y(n166),
	.B(n152),
	.A(n159), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U178 (
	.Y(n156),
	.B(n141),
	.A(n157), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U179 (
	.Y(n140),
	.B(n142),
	.A(n141), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U180 (
	.Y(n155),
	.B(i_w_full),
	.AN(i_w_inc), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U181 (
	.Y(n144),
	.B(n348),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U182 (
	.Y(n159),
	.B(n348),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U184 (
	.Y(n167),
	.B1(n340),
	.B0(n140),
	.A1N(n140),
	.A0N(\mem[15][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U185 (
	.Y(n168),
	.B1(n341),
	.B0(n140),
	.A1N(n140),
	.A0N(\mem[15][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U186 (
	.Y(n169),
	.B1(n342),
	.B0(n140),
	.A1N(n140),
	.A0N(\mem[15][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U187 (
	.Y(n170),
	.B1(n343),
	.B0(n140),
	.A1N(n140),
	.A0N(\mem[15][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U188 (
	.Y(n171),
	.B1(n344),
	.B0(n140),
	.A1N(n140),
	.A0N(\mem[15][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U189 (
	.Y(n172),
	.B1(n345),
	.B0(n140),
	.A1N(n140),
	.A0N(\mem[15][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U190 (
	.Y(n173),
	.B1(n346),
	.B0(n140),
	.A1N(n140),
	.A0N(\mem[15][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U191 (
	.Y(n174),
	.B1(n347),
	.B0(n140),
	.A1N(n140),
	.A0N(\mem[15][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U192 (
	.Y(n199),
	.B1(n148),
	.B0(n340),
	.A1N(n148),
	.A0N(\mem[11][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U193 (
	.Y(n200),
	.B1(n148),
	.B0(n341),
	.A1N(n148),
	.A0N(\mem[11][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U194 (
	.Y(n201),
	.B1(n148),
	.B0(n342),
	.A1N(n148),
	.A0N(\mem[11][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U195 (
	.Y(n202),
	.B1(n148),
	.B0(n343),
	.A1N(n148),
	.A0N(\mem[11][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U196 (
	.Y(n203),
	.B1(n148),
	.B0(n344),
	.A1N(n148),
	.A0N(\mem[11][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U197 (
	.Y(n204),
	.B1(n148),
	.B0(n345),
	.A1N(n148),
	.A0N(\mem[11][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U198 (
	.Y(n205),
	.B1(n148),
	.B0(n346),
	.A1N(n148),
	.A0N(\mem[11][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U199 (
	.Y(n206),
	.B1(n148),
	.B0(n347),
	.A1N(n148),
	.A0N(\mem[11][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U200 (
	.Y(n207),
	.B1(n150),
	.B0(n340),
	.A1N(n150),
	.A0N(\mem[10][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U201 (
	.Y(n208),
	.B1(n150),
	.B0(n341),
	.A1N(n150),
	.A0N(\mem[10][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U202 (
	.Y(n209),
	.B1(n150),
	.B0(n342),
	.A1N(n150),
	.A0N(\mem[10][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U203 (
	.Y(n210),
	.B1(n150),
	.B0(n343),
	.A1N(n150),
	.A0N(\mem[10][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U204 (
	.Y(n211),
	.B1(n150),
	.B0(n344),
	.A1N(n150),
	.A0N(\mem[10][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U205 (
	.Y(n212),
	.B1(n150),
	.B0(n345),
	.A1N(n150),
	.A0N(\mem[10][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U206 (
	.Y(n213),
	.B1(n150),
	.B0(n346),
	.A1N(n150),
	.A0N(\mem[10][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U207 (
	.Y(n214),
	.B1(n150),
	.B0(n347),
	.A1N(n150),
	.A0N(\mem[10][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U208 (
	.Y(n215),
	.B1(n151),
	.B0(n340),
	.A1N(n151),
	.A0N(\mem[9][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U209 (
	.Y(n216),
	.B1(n151),
	.B0(n341),
	.A1N(n151),
	.A0N(\mem[9][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U210 (
	.Y(n217),
	.B1(n151),
	.B0(n342),
	.A1N(n151),
	.A0N(\mem[9][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U211 (
	.Y(n218),
	.B1(n151),
	.B0(n343),
	.A1N(n151),
	.A0N(\mem[9][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U212 (
	.Y(n219),
	.B1(n151),
	.B0(n344),
	.A1N(n151),
	.A0N(\mem[9][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U213 (
	.Y(n220),
	.B1(n151),
	.B0(n345),
	.A1N(n151),
	.A0N(\mem[9][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U214 (
	.Y(n221),
	.B1(n151),
	.B0(n346),
	.A1N(n151),
	.A0N(\mem[9][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U215 (
	.Y(n222),
	.B1(n151),
	.B0(n347),
	.A1N(n151),
	.A0N(\mem[9][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U216 (
	.Y(n223),
	.B1(n154),
	.B0(n340),
	.A1N(n154),
	.A0N(\mem[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U217 (
	.Y(n224),
	.B1(n154),
	.B0(n341),
	.A1N(n154),
	.A0N(\mem[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U218 (
	.Y(n225),
	.B1(n154),
	.B0(n342),
	.A1N(n154),
	.A0N(\mem[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U219 (
	.Y(n226),
	.B1(n154),
	.B0(n343),
	.A1N(n154),
	.A0N(\mem[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U220 (
	.Y(n227),
	.B1(n154),
	.B0(n344),
	.A1N(n154),
	.A0N(\mem[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U221 (
	.Y(n228),
	.B1(n154),
	.B0(n345),
	.A1N(n154),
	.A0N(\mem[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U222 (
	.Y(n229),
	.B1(n154),
	.B0(n346),
	.A1N(n154),
	.A0N(\mem[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U223 (
	.Y(n230),
	.B1(n154),
	.B0(n347),
	.A1N(n154),
	.A0N(\mem[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U224 (
	.Y(n183),
	.B1(n145),
	.B0(n340),
	.A1N(n145),
	.A0N(\mem[13][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U225 (
	.Y(n184),
	.B1(n145),
	.B0(n341),
	.A1N(n145),
	.A0N(\mem[13][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U226 (
	.Y(n185),
	.B1(n145),
	.B0(n342),
	.A1N(n145),
	.A0N(\mem[13][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U227 (
	.Y(n186),
	.B1(n145),
	.B0(n343),
	.A1N(n145),
	.A0N(\mem[13][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U228 (
	.Y(n187),
	.B1(n145),
	.B0(n344),
	.A1N(n145),
	.A0N(\mem[13][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U229 (
	.Y(n188),
	.B1(n145),
	.B0(n345),
	.A1N(n145),
	.A0N(\mem[13][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U230 (
	.Y(n189),
	.B1(n145),
	.B0(n346),
	.A1N(n145),
	.A0N(\mem[13][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U231 (
	.Y(n190),
	.B1(n145),
	.B0(n347),
	.A1N(n145),
	.A0N(\mem[13][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U232 (
	.Y(n191),
	.B1(n147),
	.B0(n340),
	.A1N(n147),
	.A0N(\mem[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U233 (
	.Y(n192),
	.B1(n147),
	.B0(n341),
	.A1N(n147),
	.A0N(\mem[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U234 (
	.Y(n193),
	.B1(n147),
	.B0(n342),
	.A1N(n147),
	.A0N(\mem[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U235 (
	.Y(n194),
	.B1(n147),
	.B0(n343),
	.A1N(n147),
	.A0N(\mem[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U236 (
	.Y(n195),
	.B1(n147),
	.B0(n344),
	.A1N(n147),
	.A0N(\mem[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U237 (
	.Y(n196),
	.B1(n147),
	.B0(n345),
	.A1N(n147),
	.A0N(\mem[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U238 (
	.Y(n197),
	.B1(n147),
	.B0(n346),
	.A1N(n147),
	.A0N(\mem[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U239 (
	.Y(n198),
	.B1(n147),
	.B0(n347),
	.A1N(n147),
	.A0N(\mem[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U240 (
	.Y(n263),
	.B1(n162),
	.B0(n340),
	.A1N(n162),
	.A0N(\mem[3][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U241 (
	.Y(n264),
	.B1(n162),
	.B0(n341),
	.A1N(n162),
	.A0N(\mem[3][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U242 (
	.Y(n265),
	.B1(n162),
	.B0(n342),
	.A1N(n162),
	.A0N(\mem[3][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U243 (
	.Y(n266),
	.B1(n162),
	.B0(n343),
	.A1N(n162),
	.A0N(\mem[3][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U244 (
	.Y(n267),
	.B1(n162),
	.B0(n344),
	.A1N(n162),
	.A0N(\mem[3][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U245 (
	.Y(n268),
	.B1(n162),
	.B0(n345),
	.A1N(n162),
	.A0N(\mem[3][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U246 (
	.Y(n269),
	.B1(n162),
	.B0(n346),
	.A1N(n162),
	.A0N(\mem[3][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U247 (
	.Y(n270),
	.B1(n162),
	.B0(n347),
	.A1N(n162),
	.A0N(\mem[3][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U248 (
	.Y(n271),
	.B1(n163),
	.B0(n340),
	.A1N(n163),
	.A0N(\mem[2][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U249 (
	.Y(n272),
	.B1(n163),
	.B0(n341),
	.A1N(n163),
	.A0N(\mem[2][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U250 (
	.Y(n273),
	.B1(n163),
	.B0(n342),
	.A1N(n163),
	.A0N(\mem[2][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U251 (
	.Y(n274),
	.B1(n163),
	.B0(n343),
	.A1N(n163),
	.A0N(\mem[2][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U252 (
	.Y(n275),
	.B1(n163),
	.B0(n344),
	.A1N(n163),
	.A0N(\mem[2][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U253 (
	.Y(n276),
	.B1(n163),
	.B0(n345),
	.A1N(n163),
	.A0N(\mem[2][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U254 (
	.Y(n277),
	.B1(n163),
	.B0(n346),
	.A1N(n163),
	.A0N(\mem[2][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U255 (
	.Y(n278),
	.B1(n163),
	.B0(n347),
	.A1N(n163),
	.A0N(\mem[2][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U256 (
	.Y(n279),
	.B1(n164),
	.B0(n340),
	.A1N(n164),
	.A0N(\mem[1][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U257 (
	.Y(n280),
	.B1(n164),
	.B0(n341),
	.A1N(n164),
	.A0N(\mem[1][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U258 (
	.Y(n281),
	.B1(n164),
	.B0(n342),
	.A1N(n164),
	.A0N(\mem[1][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U259 (
	.Y(n282),
	.B1(n164),
	.B0(n343),
	.A1N(n164),
	.A0N(\mem[1][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U260 (
	.Y(n283),
	.B1(n164),
	.B0(n344),
	.A1N(n164),
	.A0N(\mem[1][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U261 (
	.Y(n284),
	.B1(n164),
	.B0(n345),
	.A1N(n164),
	.A0N(\mem[1][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U262 (
	.Y(n285),
	.B1(n164),
	.B0(n346),
	.A1N(n164),
	.A0N(\mem[1][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U263 (
	.Y(n286),
	.B1(n164),
	.B0(n347),
	.A1N(n164),
	.A0N(\mem[1][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U264 (
	.Y(n287),
	.B1(n166),
	.B0(n340),
	.A1N(n166),
	.A0N(\mem[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U265 (
	.Y(n288),
	.B1(n166),
	.B0(n341),
	.A1N(n166),
	.A0N(\mem[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U266 (
	.Y(n289),
	.B1(n166),
	.B0(n342),
	.A1N(n166),
	.A0N(\mem[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U267 (
	.Y(n290),
	.B1(n166),
	.B0(n343),
	.A1N(n166),
	.A0N(\mem[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U268 (
	.Y(n291),
	.B1(n166),
	.B0(n344),
	.A1N(n166),
	.A0N(\mem[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U269 (
	.Y(n292),
	.B1(n166),
	.B0(n345),
	.A1N(n166),
	.A0N(\mem[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U270 (
	.Y(n293),
	.B1(n166),
	.B0(n346),
	.A1N(n166),
	.A0N(\mem[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U271 (
	.Y(n294),
	.B1(n166),
	.B0(n347),
	.A1N(n166),
	.A0N(\mem[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U272 (
	.Y(n175),
	.B1(n143),
	.B0(n340),
	.A1N(n143),
	.A0N(\mem[14][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U273 (
	.Y(n176),
	.B1(n143),
	.B0(n341),
	.A1N(n143),
	.A0N(\mem[14][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U274 (
	.Y(n177),
	.B1(n143),
	.B0(n342),
	.A1N(n143),
	.A0N(\mem[14][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U275 (
	.Y(n178),
	.B1(n143),
	.B0(n343),
	.A1N(n143),
	.A0N(\mem[14][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U276 (
	.Y(n179),
	.B1(n143),
	.B0(n344),
	.A1N(n143),
	.A0N(\mem[14][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U277 (
	.Y(n180),
	.B1(n143),
	.B0(n345),
	.A1N(n143),
	.A0N(\mem[14][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U278 (
	.Y(n181),
	.B1(n143),
	.B0(n346),
	.A1N(n143),
	.A0N(\mem[14][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U279 (
	.Y(n182),
	.B1(n143),
	.B0(n347),
	.A1N(n143),
	.A0N(\mem[14][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U280 (
	.Y(n231),
	.B1(n156),
	.B0(n340),
	.A1N(n156),
	.A0N(\mem[7][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U281 (
	.Y(n232),
	.B1(n156),
	.B0(n341),
	.A1N(n156),
	.A0N(\mem[7][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U282 (
	.Y(n233),
	.B1(n156),
	.B0(n342),
	.A1N(n156),
	.A0N(\mem[7][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U283 (
	.Y(n234),
	.B1(n156),
	.B0(n343),
	.A1N(n156),
	.A0N(\mem[7][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U284 (
	.Y(n235),
	.B1(n156),
	.B0(n344),
	.A1N(n156),
	.A0N(\mem[7][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U285 (
	.Y(n236),
	.B1(n156),
	.B0(n345),
	.A1N(n156),
	.A0N(\mem[7][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U286 (
	.Y(n237),
	.B1(n156),
	.B0(n346),
	.A1N(n156),
	.A0N(\mem[7][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U287 (
	.Y(n238),
	.B1(n156),
	.B0(n347),
	.A1N(n156),
	.A0N(\mem[7][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U288 (
	.Y(n239),
	.B1(n158),
	.B0(n340),
	.A1N(n158),
	.A0N(\mem[6][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U289 (
	.Y(n240),
	.B1(n158),
	.B0(n341),
	.A1N(n158),
	.A0N(\mem[6][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U290 (
	.Y(n241),
	.B1(n158),
	.B0(n342),
	.A1N(n158),
	.A0N(\mem[6][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U291 (
	.Y(n242),
	.B1(n158),
	.B0(n343),
	.A1N(n158),
	.A0N(\mem[6][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U292 (
	.Y(n243),
	.B1(n158),
	.B0(n344),
	.A1N(n158),
	.A0N(\mem[6][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U293 (
	.Y(n244),
	.B1(n158),
	.B0(n345),
	.A1N(n158),
	.A0N(\mem[6][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U294 (
	.Y(n245),
	.B1(n158),
	.B0(n346),
	.A1N(n158),
	.A0N(\mem[6][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U295 (
	.Y(n246),
	.B1(n158),
	.B0(n347),
	.A1N(n158),
	.A0N(\mem[6][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U296 (
	.Y(n247),
	.B1(n160),
	.B0(n340),
	.A1N(n160),
	.A0N(\mem[5][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U297 (
	.Y(n248),
	.B1(n160),
	.B0(n341),
	.A1N(n160),
	.A0N(\mem[5][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U298 (
	.Y(n249),
	.B1(n160),
	.B0(n342),
	.A1N(n160),
	.A0N(\mem[5][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U299 (
	.Y(n250),
	.B1(n160),
	.B0(n343),
	.A1N(n160),
	.A0N(\mem[5][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U300 (
	.Y(n251),
	.B1(n160),
	.B0(n344),
	.A1N(n160),
	.A0N(\mem[5][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U301 (
	.Y(n252),
	.B1(n160),
	.B0(n345),
	.A1N(n160),
	.A0N(\mem[5][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U302 (
	.Y(n253),
	.B1(n160),
	.B0(n346),
	.A1N(n160),
	.A0N(\mem[5][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U303 (
	.Y(n254),
	.B1(n160),
	.B0(n347),
	.A1N(n160),
	.A0N(\mem[5][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U304 (
	.Y(n255),
	.B1(n161),
	.B0(n340),
	.A1N(n161),
	.A0N(\mem[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U305 (
	.Y(n256),
	.B1(n161),
	.B0(n341),
	.A1N(n161),
	.A0N(\mem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U306 (
	.Y(n257),
	.B1(n161),
	.B0(n342),
	.A1N(n161),
	.A0N(\mem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U307 (
	.Y(n258),
	.B1(n161),
	.B0(n343),
	.A1N(n161),
	.A0N(\mem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U308 (
	.Y(n259),
	.B1(n161),
	.B0(n344),
	.A1N(n161),
	.A0N(\mem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U309 (
	.Y(n260),
	.B1(n161),
	.B0(n345),
	.A1N(n161),
	.A0N(\mem[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U310 (
	.Y(n261),
	.B1(n161),
	.B0(n346),
	.A1N(n161),
	.A0N(\mem[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U311 (
	.Y(n262),
	.B1(n161),
	.B0(n347),
	.A1N(n161),
	.A0N(\mem[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U312 (
	.Y(n142),
	.B(i_wr_addr[0]),
	.A(n153), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U313 (
	.Y(n165),
	.B(i_wr_addr[3]),
	.AN(n155), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U314 (
	.Y(n157),
	.B(i_wr_addr[0]),
	.A(n165), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U315 (
	.Y(n153),
	.B(n155),
	.A(i_wr_addr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U316 (
	.Y(o_rd_data[0]),
	.S1(N12),
	.S0(N13),
	.D(n129),
	.C(n131),
	.B(n130),
	.A(n132), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U317 (
	.Y(n132),
	.S1(N11),
	.S0(N10),
	.D(\mem[3][0] ),
	.C(\mem[2][0] ),
	.B(\mem[1][0] ),
	.A(\mem[0][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U318 (
	.Y(n130),
	.S1(n318),
	.S0(N10),
	.D(\mem[11][0] ),
	.C(\mem[10][0] ),
	.B(\mem[9][0] ),
	.A(\mem[8][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U319 (
	.Y(n131),
	.S1(n318),
	.S0(N10),
	.D(\mem[7][0] ),
	.C(\mem[6][0] ),
	.B(\mem[5][0] ),
	.A(\mem[4][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U320 (
	.Y(o_rd_data[1]),
	.S1(N12),
	.S0(N13),
	.D(n133),
	.C(n135),
	.B(n134),
	.A(n136), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U321 (
	.Y(n134),
	.S1(N11),
	.S0(N10),
	.D(\mem[11][1] ),
	.C(\mem[10][1] ),
	.B(\mem[9][1] ),
	.A(\mem[8][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U322 (
	.Y(n133),
	.S1(n318),
	.S0(n321),
	.D(\mem[15][1] ),
	.C(\mem[14][1] ),
	.B(\mem[13][1] ),
	.A(\mem[12][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U323 (
	.Y(n136),
	.S1(N11),
	.S0(n321),
	.D(\mem[3][1] ),
	.C(\mem[2][1] ),
	.B(\mem[1][1] ),
	.A(\mem[0][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U324 (
	.Y(o_rd_data[2]),
	.S1(N12),
	.S0(N13),
	.D(n137),
	.C(n139),
	.B(n138),
	.A(n295), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U325 (
	.Y(n295),
	.S1(n318),
	.S0(n321),
	.D(\mem[3][2] ),
	.C(\mem[2][2] ),
	.B(\mem[1][2] ),
	.A(\mem[0][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U326 (
	.Y(n138),
	.S1(n318),
	.S0(n321),
	.D(\mem[11][2] ),
	.C(\mem[10][2] ),
	.B(\mem[9][2] ),
	.A(\mem[8][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U327 (
	.Y(n139),
	.S1(n318),
	.S0(n321),
	.D(\mem[7][2] ),
	.C(\mem[6][2] ),
	.B(\mem[5][2] ),
	.A(\mem[4][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U328 (
	.Y(o_rd_data[3]),
	.S1(N12),
	.S0(N13),
	.D(n296),
	.C(n298),
	.B(n297),
	.A(n299), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U329 (
	.Y(n299),
	.S1(n318),
	.S0(n321),
	.D(\mem[3][3] ),
	.C(\mem[2][3] ),
	.B(\mem[1][3] ),
	.A(\mem[0][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U330 (
	.Y(n297),
	.S1(n318),
	.S0(n321),
	.D(\mem[11][3] ),
	.C(\mem[10][3] ),
	.B(\mem[9][3] ),
	.A(\mem[8][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U331 (
	.Y(n298),
	.S1(n318),
	.S0(n321),
	.D(\mem[7][3] ),
	.C(\mem[6][3] ),
	.B(\mem[5][3] ),
	.A(\mem[4][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U332 (
	.Y(o_rd_data[4]),
	.S1(N12),
	.S0(N13),
	.D(n300),
	.C(n302),
	.B(n301),
	.A(n303), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U333 (
	.Y(n303),
	.S1(n318),
	.S0(n322),
	.D(\mem[3][4] ),
	.C(\mem[2][4] ),
	.B(\mem[1][4] ),
	.A(\mem[0][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U334 (
	.Y(n301),
	.S1(n318),
	.S0(n321),
	.D(\mem[11][4] ),
	.C(\mem[10][4] ),
	.B(\mem[9][4] ),
	.A(\mem[8][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U335 (
	.Y(n302),
	.S1(n318),
	.S0(n321),
	.D(\mem[7][4] ),
	.C(\mem[6][4] ),
	.B(\mem[5][4] ),
	.A(\mem[4][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U336 (
	.Y(o_rd_data[5]),
	.S1(N12),
	.S0(N13),
	.D(n304),
	.C(n306),
	.B(n305),
	.A(n307), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U337 (
	.Y(n307),
	.S1(N11),
	.S0(n322),
	.D(\mem[3][5] ),
	.C(\mem[2][5] ),
	.B(\mem[1][5] ),
	.A(\mem[0][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U338 (
	.Y(n305),
	.S1(N11),
	.S0(n322),
	.D(\mem[11][5] ),
	.C(\mem[10][5] ),
	.B(\mem[9][5] ),
	.A(\mem[8][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U339 (
	.Y(n306),
	.S1(N11),
	.S0(n322),
	.D(\mem[7][5] ),
	.C(\mem[6][5] ),
	.B(\mem[5][5] ),
	.A(\mem[4][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U340 (
	.Y(o_rd_data[6]),
	.S1(N12),
	.S0(N13),
	.D(n308),
	.C(n310),
	.B(n309),
	.A(n311), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U341 (
	.Y(n311),
	.S1(N11),
	.S0(n322),
	.D(\mem[3][6] ),
	.C(\mem[2][6] ),
	.B(\mem[1][6] ),
	.A(\mem[0][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U342 (
	.Y(n309),
	.S1(N11),
	.S0(n322),
	.D(\mem[11][6] ),
	.C(\mem[10][6] ),
	.B(\mem[9][6] ),
	.A(\mem[8][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U343 (
	.Y(n310),
	.S1(N11),
	.S0(n322),
	.D(\mem[7][6] ),
	.C(\mem[6][6] ),
	.B(\mem[5][6] ),
	.A(\mem[4][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U344 (
	.Y(o_rd_data[7]),
	.S1(N12),
	.S0(N13),
	.D(n312),
	.C(n314),
	.B(n313),
	.A(n315), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U345 (
	.Y(n315),
	.S1(N11),
	.S0(n322),
	.D(\mem[3][7] ),
	.C(\mem[2][7] ),
	.B(\mem[1][7] ),
	.A(\mem[0][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U346 (
	.Y(n313),
	.S1(N11),
	.S0(n322),
	.D(\mem[11][7] ),
	.C(\mem[10][7] ),
	.B(\mem[9][7] ),
	.A(\mem[8][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U347 (
	.Y(n314),
	.S1(N11),
	.S0(n322),
	.D(\mem[7][7] ),
	.C(\mem[6][7] ),
	.B(\mem[5][7] ),
	.A(\mem[4][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U348 (
	.Y(n135),
	.S1(n318),
	.S0(n321),
	.D(\mem[7][1] ),
	.C(\mem[6][1] ),
	.B(\mem[5][1] ),
	.A(\mem[4][1] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U349 (
	.Y(n129),
	.S1(n318),
	.S0(n322),
	.D(\mem[15][0] ),
	.C(\mem[14][0] ),
	.B(\mem[13][0] ),
	.A(\mem[12][0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U350 (
	.Y(n137),
	.S1(n318),
	.S0(n321),
	.D(\mem[15][2] ),
	.C(\mem[14][2] ),
	.B(\mem[13][2] ),
	.A(\mem[12][2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U351 (
	.Y(n296),
	.S1(n318),
	.S0(n321),
	.D(\mem[15][3] ),
	.C(\mem[14][3] ),
	.B(\mem[13][3] ),
	.A(\mem[12][3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U352 (
	.Y(n300),
	.S1(n318),
	.S0(n321),
	.D(\mem[15][4] ),
	.C(\mem[14][4] ),
	.B(\mem[13][4] ),
	.A(\mem[12][4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U353 (
	.Y(n304),
	.S1(N11),
	.S0(n322),
	.D(\mem[15][5] ),
	.C(\mem[14][5] ),
	.B(\mem[13][5] ),
	.A(\mem[12][5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U354 (
	.Y(n308),
	.S1(N11),
	.S0(n322),
	.D(\mem[15][6] ),
	.C(\mem[14][6] ),
	.B(\mem[13][6] ),
	.A(\mem[12][6] ), 
	.VDD(VDD), 
	.VSS(VSS));
   MX4X1M U355 (
	.Y(n312),
	.S1(N11),
	.S0(n322),
	.D(\mem[15][7] ),
	.C(\mem[14][7] ),
	.B(\mem[13][7] ),
	.A(\mem[12][7] ), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U356 (
	.Y(n316),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U357 (
	.Y(n350),
	.A(i_wr_addr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U358 (
	.Y(n349),
	.A(i_wr_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U359 (
	.Y(n348),
	.A(i_wr_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U360 (
	.Y(n354),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U361 (
	.Y(n355),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U362 (
	.Y(n356),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   DLY1X4M U363 (
	.Y(n357),
	.A(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_ADDR_WIDTH4_test_1 (
	i_clk, 
	i_rst_n, 
	i_r_d_ptr, 
	wq2_r_d_ptr, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input i_clk;
   input i_rst_n;
   input [4:0] i_r_d_ptr;
   output [4:0] wq2_r_d_ptr;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [4:0] R1;

   // Module instantiations
   SDFFRQX2M \R2_reg[2]  (
	.SI(wq2_r_d_ptr[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[2]),
	.D(R1[2]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R2_reg[0]  (
	.SI(R1[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[0]),
	.D(R1[0]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R2_reg[1]  (
	.SI(wq2_r_d_ptr[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[1]),
	.D(R1[1]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R2_reg[4]  (
	.SI(wq2_r_d_ptr[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[4]),
	.D(R1[4]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R2_reg[3]  (
	.SI(wq2_r_d_ptr[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[3]),
	.D(R1[3]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[4]  (
	.SI(R1[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[4]),
	.D(i_r_d_ptr[4]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[3]  (
	.SI(R1[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[3]),
	.D(i_r_d_ptr[3]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[2]  (
	.SI(R1[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[2]),
	.D(i_r_d_ptr[2]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[1]  (
	.SI(R1[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[1]),
	.D(i_r_d_ptr[1]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[0]),
	.D(i_r_d_ptr[0]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DF_SYNC_ADDR_WIDTH4_test_0 (
	i_clk, 
	i_rst_n, 
	i_r_d_ptr, 
	wq2_r_d_ptr, 
	test_si, 
	test_se, 
	CLK_R_M__L5_N4, 
	VDD, 
	VSS);
   input i_clk;
   input i_rst_n;
   input [4:0] i_r_d_ptr;
   output [4:0] wq2_r_d_ptr;
   input test_si;
   input test_se;
   input CLK_R_M__L5_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire [4:0] R1;

   // Module instantiations
   SDFFRQX2M \R2_reg[4]  (
	.SI(wq2_r_d_ptr[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[4]),
	.D(R1[4]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R2_reg[3]  (
	.SI(wq2_r_d_ptr[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[3]),
	.D(R1[3]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R2_reg[2]  (
	.SI(wq2_r_d_ptr[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[2]),
	.D(R1[2]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R2_reg[1]  (
	.SI(wq2_r_d_ptr[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[1]),
	.D(R1[1]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R2_reg[0]  (
	.SI(R1[4]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(wq2_r_d_ptr[0]),
	.D(R1[0]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[4]  (
	.SI(R1[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[4]),
	.D(i_r_d_ptr[4]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[3]  (
	.SI(R1[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[3]),
	.D(i_r_d_ptr[3]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[2]  (
	.SI(R1[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[2]),
	.D(i_r_d_ptr[2]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[1]  (
	.SI(R1[0]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[1]),
	.D(i_r_d_ptr[1]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \R1_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(R1[0]),
	.D(i_r_d_ptr[0]),
	.CK(i_clk), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_RD_DATA_WIDTH8_ADDR_WIDTH4_test_1 (
	i_r_clk, 
	i_rst_n, 
	i_r_inc, 
	rq2_wptr, 
	o_r_empty, 
	o_rd_addr, 
	o_rptr, 
	test_si2, 
	test_si1, 
	test_se, 
	TX_CLK_M__L3_N1, 
	VDD, 
	VSS);
   input i_r_clk;
   input i_rst_n;
   input i_r_inc;
   input [4:0] rq2_wptr;
   output o_r_empty;
   output [3:0] o_rd_addr;
   output [4:0] o_rptr;
   input test_si2;
   input test_si1;
   input test_se;
   input TX_CLK_M__L3_N1;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire n1;
   wire n3;
   wire n5;
   wire n7;
   wire n9;
   wire n11;
   wire \add_23/carry[4] ;
   wire \add_23/carry[3] ;
   wire \add_23/carry[2] ;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;

   // Module instantiations
   SDFFRQX2M \o_rptr_reg_reg[4]  (
	.SI(o_rd_addr[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(o_rptr[4]),
	.D(n9),
	.CK(i_r_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \o_rptr_reg_reg[0]  (
	.SI(test_si1),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(o_rd_addr[0]),
	.D(n11),
	.CK(i_r_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \o_rptr_reg_reg[1]  (
	.SI(test_si2),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(o_rd_addr[1]),
	.D(n7),
	.CK(TX_CLK_M__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \o_rptr_reg_reg[2]  (
	.SI(o_rd_addr[1]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(o_rd_addr[2]),
	.D(n5),
	.CK(TX_CLK_M__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \o_rptr_reg_reg[3]  (
	.SI(o_rd_addr[2]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(o_rd_addr[3]),
	.D(n3),
	.CK(TX_CLK_M__L3_N1), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U3 (
	.Y(n11),
	.B1(n1),
	.B0(n12),
	.A1N(n1),
	.A0(o_rd_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U4 (
	.Y(n1),
	.B(o_r_empty),
	.AN(i_r_inc), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U5 (
	.Y(n3),
	.B1(n1),
	.B0(N6),
	.A1N(n1),
	.A0(o_rd_addr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U6 (
	.Y(n5),
	.B1(n1),
	.B0(N5),
	.A1N(n1),
	.A0(o_rd_addr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U7 (
	.Y(n7),
	.B1(n1),
	.B0(N4),
	.A1N(n1),
	.A0(o_rd_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U8 (
	.Y(n9),
	.B1(n1),
	.B0(N7),
	.A1N(n1),
	.A0(o_rptr[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n12),
	.A(o_rd_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U10 (
	.Y(o_rptr[2]),
	.B(o_rd_addr[2]),
	.A(o_rd_addr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U11 (
	.Y(o_rptr[1]),
	.B(o_rd_addr[1]),
	.A(o_rd_addr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U12 (
	.Y(o_rptr[0]),
	.B(o_rd_addr[0]),
	.A(o_rd_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U18 (
	.Y(o_rptr[3]),
	.B(o_rd_addr[3]),
	.A(o_rptr[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U19 (
	.S(N5),
	.CO(\add_23/carry[3] ),
	.B(\add_23/carry[2] ),
	.A(o_rd_addr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U20 (
	.S(N4),
	.CO(\add_23/carry[2] ),
	.B(o_rd_addr[0]),
	.A(o_rd_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U21 (
	.S(N6),
	.CO(\add_23/carry[4] ),
	.B(\add_23/carry[3] ),
	.A(o_rd_addr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(N7),
	.B(o_rptr[4]),
	.A(\add_23/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(n20),
	.B(o_rptr[2]),
	.A(rq2_wptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U24 (
	.Y(n13),
	.B(o_rptr[0]),
	.AN(rq2_wptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U25 (
	.Y(n16),
	.B1(n13),
	.B0(rq2_wptr[1]),
	.A1N(o_rptr[1]),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U26 (
	.Y(n14),
	.B(rq2_wptr[0]),
	.AN(o_rptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U27 (
	.Y(n15),
	.B1(n14),
	.B0(o_rptr[1]),
	.A1N(rq2_wptr[1]),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U28 (
	.Y(n19),
	.B(n15),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U29 (
	.Y(n18),
	.B(o_rptr[3]),
	.A(rq2_wptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U30 (
	.Y(n17),
	.B(o_rptr[4]),
	.A(rq2_wptr[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U31 (
	.Y(o_r_empty),
	.D(n17),
	.C(n18),
	.B(n19),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FIFO_WR_DATA_WIDTH8_ADDR_WIDTH4_test_1 (
	i_w_clk, 
	i_rst_n, 
	i_w_inc, 
	wq2_rptr, 
	o_w_full, 
	o_wr_addr, 
	o_wptr, 
	test_si, 
	test_se, 
	FE_OFN2_RST_SYNC_1_mux, 
	CLK_R_M__L5_N3, 
	VDD, 
	VSS);
   input i_w_clk;
   input i_rst_n;
   input i_w_inc;
   input [4:0] wq2_rptr;
   output o_w_full;
   output [3:0] o_wr_addr;
   output [4:0] o_wptr;
   input test_si;
   input test_se;
   input FE_OFN2_RST_SYNC_1_mux;
   input CLK_R_M__L5_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N3;
   wire N4;
   wire N5;
   wire N6;
   wire N7;
   wire n7;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire \add_22/carry[4] ;
   wire \add_22/carry[3] ;
   wire \add_22/carry[2] ;
   wire n8;
   wire n21;

   // Module instantiations
   SDFFRQX2M \o_wptr_reg_reg[4]  (
	.SI(o_wr_addr[3]),
	.SE(test_se),
	.RN(i_rst_n),
	.Q(o_wptr[4]),
	.D(n19),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \o_wptr_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(o_wr_addr[0]),
	.D(n20),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \o_wptr_reg_reg[3]  (
	.SI(o_wr_addr[2]),
	.SE(test_se),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(o_wr_addr[3]),
	.D(n16),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \o_wptr_reg_reg[1]  (
	.SI(N3),
	.SE(test_se),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.Q(o_wr_addr[1]),
	.D(n18),
	.CK(i_w_clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRX1M \o_wptr_reg_reg[2]  (
	.SI(o_wr_addr[1]),
	.SE(test_se),
	.RN(FE_OFN2_RST_SYNC_1_mux),
	.QN(n7),
	.Q(o_wr_addr[2]),
	.D(n17),
	.CK(CLK_R_M__L5_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U9 (
	.Y(n9),
	.B(o_w_full),
	.AN(i_w_inc), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U10 (
	.Y(n16),
	.B1(n21),
	.B0(n9),
	.A1N(n9),
	.A0N(N6), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U11 (
	.Y(n18),
	.B1(n8),
	.B0(n9),
	.A1N(n9),
	.A0N(N4), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U12 (
	.Y(o_w_full),
	.D(n13),
	.C(n12),
	.B(n11),
	.A(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U13 (
	.Y(n11),
	.B(wq2_rptr[1]),
	.A(o_wptr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U14 (
	.Y(n10),
	.B(wq2_rptr[0]),
	.A(o_wptr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U15 (
	.Y(n13),
	.B(wq2_rptr[2]),
	.A(o_wptr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n8),
	.A(o_wr_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n21),
	.A(o_wr_addr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U18 (
	.Y(n12),
	.B(n15),
	.A(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U19 (
	.Y(n15),
	.B(wq2_rptr[4]),
	.A(o_wptr[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U20 (
	.Y(n14),
	.B(wq2_rptr[3]),
	.A(o_wptr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U21 (
	.Y(o_wptr[0]),
	.B(o_wr_addr[1]),
	.A(o_wr_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(o_wptr[1]),
	.B(n7),
	.A(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(o_wptr[3]),
	.B(o_wr_addr[3]),
	.A(o_wptr[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U24 (
	.Y(o_wptr[2]),
	.B(n21),
	.A(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U25 (
	.Y(n17),
	.B1(n7),
	.B0(n9),
	.A1N(n9),
	.A0N(N5), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U26 (
	.Y(n19),
	.B1(n9),
	.B0(N7),
	.A1N(n9),
	.A0(o_wptr[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U27 (
	.Y(n20),
	.B1(n9),
	.B0(N3),
	.A1N(n9),
	.A0(o_wr_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(N3),
	.A(o_wr_addr[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U29 (
	.S(N5),
	.CO(\add_22/carry[3] ),
	.B(\add_22/carry[2] ),
	.A(o_wr_addr[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U30 (
	.S(N4),
	.CO(\add_22/carry[2] ),
	.B(o_wr_addr[0]),
	.A(o_wr_addr[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U31 (
	.S(N6),
	.CO(\add_22/carry[4] ),
	.B(\add_22/carry[3] ),
	.A(o_wr_addr[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U32 (
	.Y(N7),
	.B(o_wptr[4]),
	.A(\add_22/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module DATA_SYNC_test_1 (
	clk, 
	rst_n, 
	unsync_bus, 
	bus_enable, 
	sync_bus, 
	enable_pulse, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input clk;
   input rst_n;
   input [7:0] unsync_bus;
   input bus_enable;
   output [7:0] sync_bus;
   output enable_pulse;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire enable_pulse_gen_reg;
   wire n1;
   wire n3;
   wire n5;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n22;
   wire [1:0] sync_reg;

   assign test_so = sync_reg[1] ;

   // Module instantiations
   SDFFRQX2M enable_pulse_gen_reg_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(rst_n),
	.Q(enable_pulse_gen_reg),
	.D(sync_reg[1]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[1]  (
	.SI(sync_reg[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_reg[1]),
	.D(sync_reg[0]),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[0]  (
	.SI(enable_pulse),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[0]),
	.D(n3),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[7]  (
	.SI(sync_bus[6]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[7]),
	.D(n17),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[6]  (
	.SI(sync_bus[5]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[6]),
	.D(n15),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[3]  (
	.SI(sync_bus[2]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[3]),
	.D(n9),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[2]  (
	.SI(sync_bus[1]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[2]),
	.D(n7),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[4]  (
	.SI(sync_bus[3]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[4]),
	.D(n11),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[5]  (
	.SI(sync_bus[4]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[5]),
	.D(n13),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_bus_reg[1]  (
	.SI(sync_bus[0]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_bus[1]),
	.D(n5),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M enable_pulse_reg (
	.SI(enable_pulse_gen_reg),
	.SE(test_se),
	.RN(rst_n),
	.Q(enable_pulse),
	.D(n22),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \sync_reg_reg[0]  (
	.SI(sync_bus[7]),
	.SE(test_se),
	.RN(rst_n),
	.Q(sync_reg[0]),
	.D(bus_enable),
	.CK(clk), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U3 (
	.Y(n22),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX2M U4 (
	.Y(n1),
	.B(sync_reg[1]),
	.AN(enable_pulse_gen_reg), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U5 (
	.Y(n3),
	.B1(n1),
	.B0(sync_bus[0]),
	.A1(n22),
	.A0(unsync_bus[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U6 (
	.Y(n5),
	.B1(n1),
	.B0(sync_bus[1]),
	.A1(n22),
	.A0(unsync_bus[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U7 (
	.Y(n7),
	.B1(n1),
	.B0(sync_bus[2]),
	.A1(n22),
	.A0(unsync_bus[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U8 (
	.Y(n9),
	.B1(n1),
	.B0(sync_bus[3]),
	.A1(n22),
	.A0(unsync_bus[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U9 (
	.Y(n11),
	.B1(n1),
	.B0(sync_bus[4]),
	.A1(n22),
	.A0(unsync_bus[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U10 (
	.Y(n13),
	.B1(n1),
	.B0(sync_bus[5]),
	.A1(n22),
	.A0(unsync_bus[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U11 (
	.Y(n15),
	.B1(n1),
	.B0(sync_bus[6]),
	.A1(n22),
	.A0(unsync_bus[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U12 (
	.Y(n17),
	.B1(n1),
	.B0(sync_bus[7]),
	.A1(n22),
	.A0(unsync_bus[7]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module RX_TOP_test_1 (
	CLK_RX, 
	RST_RX, 
	RX_IN_RX, 
	PAR_EN_RX, 
	PAR_TYP_RX, 
	prescale_RX, 
	P_DATA_RX, 
	data_valid_RX, 
	parity_error_RX, 
	stop_error_RX, 
	test_si1, 
	test_so1, 
	test_se, 
	FE_OFN4_RST_SYNC_2_mux, 
	VDD, 
	VSS);
   input CLK_RX;
   input RST_RX;
   input RX_IN_RX;
   input PAR_EN_RX;
   input PAR_TYP_RX;
   input [5:0] prescale_RX;
   output [7:0] P_DATA_RX;
   output data_valid_RX;
   output parity_error_RX;
   output stop_error_RX;
   input test_si1;
   output test_so1;
   input test_se;
   input FE_OFN4_RST_SYNC_2_mux;
   inout VDD;
   inout VSS;

   // Internal wires
   wire strt_chk_en_wire;
   wire sample_bit_wire;
   wire strt_glitch_wire;
   wire par_chk_en_wire;
   wire stp_chk_en_wire;
   wire deser_en_wire;
   wire data_samp_en_wire;
   wire enable_wire;
   wire n3;
   wire n4;
   wire [5:0] edge_cnt_wires;
   wire [5:0] bit_cnt_wires;

   assign test_so1 = strt_glitch_wire ;

   // Module instantiations
   strt_check_RX_test_1 strt_check_RX1 (
	.CLK_start(CLK_RX),
	.RST_start(RST_RX),
	.strt_chk_en(strt_chk_en_wire),
	.sample_bit_par_chk(sample_bit_wire),
	.strt_glitch_chk(strt_glitch_wire),
	.test_si(parity_error_RX),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_check_RX_test_1 parity_check_RX1 (
	.CLK_par(CLK_RX),
	.RST_par(RST_RX),
	.P_DATA_par_chk({ P_DATA_RX[7],
		P_DATA_RX[6],
		P_DATA_RX[5],
		P_DATA_RX[4],
		P_DATA_RX[3],
		P_DATA_RX[2],
		P_DATA_RX[1],
		P_DATA_RX[0] }),
	.PAR_TYP_par_chk(PAR_TYP_RX),
	.par_chk_en(par_chk_en_wire),
	.sample_bit_par_chk(sample_bit_wire),
	.par_err(parity_error_RX),
	.test_si(edge_cnt_wires[5]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   stop_check_RX_test_1 stop_check_RX1 (
	.CLK_stop(CLK_RX),
	.RST_stop(RST_RX),
	.stp_chk_en(stp_chk_en_wire),
	.sample_bit_par_chk(sample_bit_wire),
	.Stop_Error(stop_error_RX),
	.test_si(prescale_RX[0]),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   deserializer_RX_test_1 deserializer_RX1 (
	.CLK_des(CLK_RX),
	.RST_des(RST_RX),
	.sample_bit_deser(sample_bit_wire),
	.deser_en(deser_en_wire),
	.edge_cnt({ edge_cnt_wires[5],
		edge_cnt_wires[4],
		edge_cnt_wires[3],
		edge_cnt_wires[2],
		edge_cnt_wires[1],
		edge_cnt_wires[0] }),
	.prescale_FSM({ prescale_RX[5],
		prescale_RX[4],
		prescale_RX[3],
		prescale_RX[2],
		prescale_RX[1],
		prescale_RX[0] }),
	.P_DATA_des({ P_DATA_RX[7],
		P_DATA_RX[6],
		P_DATA_RX[5],
		P_DATA_RX[4],
		P_DATA_RX[3],
		P_DATA_RX[2],
		P_DATA_RX[1],
		P_DATA_RX[0] }),
	.test_so(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   data_sampling_RX_test_1 data_sampling_RX1 (
	.CLK_SAM(CLK_RX),
	.RST_SAM(RST_RX),
	.RX_IN(RX_IN_RX),
	.data_samp_en(data_samp_en_wire),
	.edge_cnt({ edge_cnt_wires[5],
		edge_cnt_wires[4],
		edge_cnt_wires[3],
		edge_cnt_wires[2],
		edge_cnt_wires[1],
		edge_cnt_wires[0] }),
	.prescale({ prescale_RX[5],
		prescale_RX[4],
		prescale_RX[3],
		prescale_RX[2],
		prescale_RX[1],
		prescale_RX[0] }),
	.sample_bit_samp(sample_bit_wire),
	.test_si(n4),
	.test_se(test_se),
	.FE_OFN4_RST_SYNC_2_mux(FE_OFN4_RST_SYNC_2_mux), 
	.VDD(VDD), 
	.VSS(VSS));
   edge_bit_counter_RX_test_1 edge_bit_counter_RX1 (
	.CLK_EDGE(CLK_RX),
	.RST_EDGE(FE_OFN4_RST_SYNC_2_mux),
	.enable_edge(enable_wire),
	.prescale_edge({ prescale_RX[5],
		prescale_RX[4],
		prescale_RX[3],
		prescale_RX[2],
		prescale_RX[1],
		prescale_RX[0] }),
	.bit_cnt_edge({ bit_cnt_wires[5],
		bit_cnt_wires[4],
		bit_cnt_wires[3],
		bit_cnt_wires[2],
		bit_cnt_wires[1],
		bit_cnt_wires[0] }),
	.edge_cnt_edge({ edge_cnt_wires[5],
		edge_cnt_wires[4],
		edge_cnt_wires[3],
		edge_cnt_wires[2],
		edge_cnt_wires[1],
		edge_cnt_wires[0] }),
	.test_si(n3),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   FSM_RX_test_1 FSM_RX1 (
	.CLK_FSM(CLK_RX),
	.RST_FSM(RST_RX),
	.RX_IN(RX_IN_RX),
	.bit_cnt_FSM({ bit_cnt_wires[5],
		bit_cnt_wires[4],
		bit_cnt_wires[3],
		bit_cnt_wires[2],
		bit_cnt_wires[1],
		bit_cnt_wires[0] }),
	.edge_cnt_FSM({ edge_cnt_wires[5],
		edge_cnt_wires[4],
		edge_cnt_wires[3],
		edge_cnt_wires[2],
		edge_cnt_wires[1],
		edge_cnt_wires[0] }),
	.PAR_EN_FSM(PAR_EN_RX),
	.par_err_FSM(parity_error_RX),
	.strt_glitch_FSM(strt_glitch_wire),
	.stp_err_FSM(stop_error_RX),
	.prescale_FSM({ prescale_RX[5],
		prescale_RX[4],
		prescale_RX[3],
		prescale_RX[2],
		prescale_RX[1],
		prescale_RX[0] }),
	.par_chk_en_FSM(par_chk_en_wire),
	.strt_chk_en_FSM(strt_chk_en_wire),
	.stp_chk_en_FSM(stp_chk_en_wire),
	.enable_FSM(enable_wire),
	.data_samp_en_FSM(data_samp_en_wire),
	.data_valid_FSM(data_valid_RX),
	.deser_en_FSM(deser_en_wire),
	.test_si(test_si1),
	.test_so(n4),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module strt_check_RX_test_1 (
	CLK_start, 
	RST_start, 
	strt_chk_en, 
	sample_bit_par_chk, 
	strt_glitch_chk, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK_start;
   input RST_start;
   input strt_chk_en;
   input sample_bit_par_chk;
   output strt_glitch_chk;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire strt_glitch_chk_reg;

   // Module instantiations
   SDFFRQX2M strt_glitch_chk_reg_inst (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_start),
	.Q(strt_glitch_chk),
	.D(strt_glitch_chk_reg),
	.CK(CLK_start), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U4 (
	.Y(strt_glitch_chk_reg),
	.B(sample_bit_par_chk),
	.A(strt_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_check_RX_test_1 (
	CLK_par, 
	RST_par, 
	P_DATA_par_chk, 
	PAR_TYP_par_chk, 
	par_chk_en, 
	sample_bit_par_chk, 
	par_err, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK_par;
   input RST_par;
   input [7:0] P_DATA_par_chk;
   input PAR_TYP_par_chk;
   input par_chk_en;
   input sample_bit_par_chk;
   output par_err;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n9;
   wire n2;

   // Module instantiations
   SDFFRQX4M par_err_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_par),
	.Q(par_err),
	.D(n9),
	.CK(CLK_par), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U2 (
	.Y(n9),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(par_err), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U3 (
	.Y(n1),
	.C(n5),
	.B(n4),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n2),
	.A(par_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U5 (
	.Y(n5),
	.B(PAR_TYP_par_chk),
	.A(sample_bit_par_chk), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U6 (
	.Y(n4),
	.C(n6),
	.B(P_DATA_par_chk[4]),
	.A(P_DATA_par_chk[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U7 (
	.Y(n6),
	.B(P_DATA_par_chk[6]),
	.A(P_DATA_par_chk[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U8 (
	.Y(n3),
	.C(n7),
	.B(P_DATA_par_chk[0]),
	.A(P_DATA_par_chk[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U9 (
	.Y(n7),
	.B(P_DATA_par_chk[2]),
	.A(P_DATA_par_chk[3]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module stop_check_RX_test_1 (
	CLK_stop, 
	RST_stop, 
	stp_chk_en, 
	sample_bit_par_chk, 
	Stop_Error, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK_stop;
   input RST_stop;
   input stp_chk_en;
   input sample_bit_par_chk;
   output Stop_Error;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire stp_err_chk;

   // Module instantiations
   SDFFRQX4M Stop_Error_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_stop),
	.Q(Stop_Error),
	.D(stp_err_chk),
	.CK(CLK_stop), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U4 (
	.Y(stp_err_chk),
	.B(sample_bit_par_chk),
	.AN(stp_chk_en), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module deserializer_RX_test_1 (
	CLK_des, 
	RST_des, 
	sample_bit_deser, 
	deser_en, 
	edge_cnt, 
	prescale_FSM, 
	P_DATA_des, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK_des;
   input RST_des;
   input sample_bit_deser;
   input deser_en;
   input [5:0] edge_cnt;
   input [5:0] prescale_FSM;
   output [7:0] P_DATA_des;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n10;
   wire n12;
   wire n14;
   wire n16;
   wire n18;
   wire n20;
   wire n22;
   wire n24;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n25;

   assign test_so = n3 ;

   // Module instantiations
   SDFFRQX2M \P_DATA_des_reg[0]  (
	.SI(sample_bit_deser),
	.SE(test_se),
	.RN(RST_des),
	.Q(P_DATA_des[0]),
	.D(n10),
	.CK(CLK_des), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_des_reg[5]  (
	.SI(n6),
	.SE(test_se),
	.RN(RST_des),
	.Q(P_DATA_des[5]),
	.D(n20),
	.CK(CLK_des), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_des_reg[1]  (
	.SI(P_DATA_des[0]),
	.SE(test_se),
	.RN(RST_des),
	.Q(P_DATA_des[1]),
	.D(n12),
	.CK(CLK_des), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_des_reg[4]  (
	.SI(n7),
	.SE(test_se),
	.RN(RST_des),
	.Q(P_DATA_des[4]),
	.D(n18),
	.CK(CLK_des), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_des_reg[7]  (
	.SI(n4),
	.SE(test_se),
	.RN(RST_des),
	.Q(P_DATA_des[7]),
	.D(n24),
	.CK(CLK_des), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_des_reg[3]  (
	.SI(n8),
	.SE(test_se),
	.RN(RST_des),
	.Q(P_DATA_des[3]),
	.D(n16),
	.CK(CLK_des), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_des_reg[6]  (
	.SI(n5),
	.SE(test_se),
	.RN(RST_des),
	.Q(P_DATA_des[6]),
	.D(n22),
	.CK(CLK_des), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \P_DATA_des_reg[2]  (
	.SI(n25),
	.SE(test_se),
	.RN(RST_des),
	.Q(P_DATA_des[2]),
	.D(n14),
	.CK(CLK_des), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U2 (
	.Y(n2),
	.A(deser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U4 (
	.Y(n12),
	.B1(n25),
	.B0(deser_en),
	.A1(n8),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U5 (
	.Y(n14),
	.B1(n8),
	.B0(deser_en),
	.A1(n7),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U6 (
	.Y(n16),
	.B1(n7),
	.B0(deser_en),
	.A1(n6),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U7 (
	.Y(n18),
	.B1(n6),
	.B0(deser_en),
	.A1(n5),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U8 (
	.Y(n20),
	.B1(n5),
	.B0(deser_en),
	.A1(n4),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U9 (
	.Y(n22),
	.B1(n4),
	.B0(deser_en),
	.A1(n3),
	.A0(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U10 (
	.Y(n10),
	.B1(n2),
	.B0(n25),
	.A1N(n2),
	.A0N(P_DATA_des[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U11 (
	.Y(n24),
	.B1(n3),
	.B0(deser_en),
	.A1N(deser_en),
	.A0N(sample_bit_deser), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n8),
	.A(P_DATA_des[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n4),
	.A(P_DATA_des[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U14 (
	.Y(n3),
	.A(P_DATA_des[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n7),
	.A(P_DATA_des[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n25),
	.A(P_DATA_des[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n6),
	.A(P_DATA_des[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n5),
	.A(P_DATA_des[5]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module data_sampling_RX_test_1 (
	CLK_SAM, 
	RST_SAM, 
	RX_IN, 
	data_samp_en, 
	edge_cnt, 
	prescale, 
	sample_bit_samp, 
	test_si, 
	test_se, 
	FE_OFN4_RST_SYNC_2_mux, 
	VDD, 
	VSS);
   input CLK_SAM;
   input RST_SAM;
   input RX_IN;
   input data_samp_en;
   input [5:0] edge_cnt;
   input [5:0] prescale;
   output sample_bit_samp;
   input test_si;
   input test_se;
   input FE_OFN4_RST_SYNC_2_mux;
   inout VDD;
   inout VSS;

   // Internal wires
   wire \RX_IN_reg[0] ;
   wire N11;
   wire N12;
   wire N13;
   wire N14;
   wire N15;
   wire N16;
   wire N18;
   wire N25;
   wire n27;
   wire n28;
   wire n29;
   wire \sub_29/carry[5] ;
   wire \sub_29/carry[4] ;
   wire \sub_29/carry[3] ;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;

   assign N11 = prescale[0] ;

   // Module instantiations
   SDFFRQX2M \RX_IN_reg_reg[1]  (
	.SI(\RX_IN_reg[0] ),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(N25),
	.D(n28),
	.CK(CLK_SAM), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \RX_IN_reg_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_SAM),
	.Q(\RX_IN_reg[0] ),
	.D(n29),
	.CK(CLK_SAM), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX1M sample_bit_samp_reg (
	.SN(FE_OFN4_RST_SYNC_2_mux),
	.SI(N25),
	.SE(test_se),
	.Q(sample_bit_samp),
	.D(n27),
	.CK(CLK_SAM), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U7 (
	.Y(n2),
	.B(\sub_29/carry[5] ),
	.A(prescale[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(N12),
	.A(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U9 (
	.Y(N16),
	.B(prescale[5]),
	.A(\sub_29/carry[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U10 (
	.Y(\sub_29/carry[5] ),
	.B(\sub_29/carry[4] ),
	.A(prescale[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U11 (
	.Y(N15),
	.B(prescale[4]),
	.A(\sub_29/carry[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U12 (
	.Y(\sub_29/carry[4] ),
	.B(\sub_29/carry[3] ),
	.A(prescale[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U13 (
	.Y(N14),
	.B(prescale[3]),
	.A(\sub_29/carry[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U14 (
	.Y(\sub_29/carry[3] ),
	.B(prescale[1]),
	.A(prescale[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U15 (
	.Y(N13),
	.B(prescale[2]),
	.A(prescale[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U16 (
	.Y(n3),
	.B(edge_cnt[0]),
	.AN(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U17 (
	.Y(n7),
	.B1(n3),
	.B0(N12),
	.A1N(edge_cnt[1]),
	.A0(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U18 (
	.Y(n6),
	.B(edge_cnt[5]),
	.A(N16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U19 (
	.Y(n4),
	.B(N11),
	.AN(edge_cnt[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U20 (
	.Y(n5),
	.B1(n4),
	.B0(edge_cnt[1]),
	.A1N(N12),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U21 (
	.Y(n11),
	.D(n5),
	.C(n6),
	.B(n7),
	.AN(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U22 (
	.Y(n10),
	.B(edge_cnt[4]),
	.A(N15), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U23 (
	.Y(n9),
	.B(edge_cnt[2]),
	.A(N13), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U24 (
	.Y(n8),
	.B(edge_cnt[3]),
	.A(N14), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U25 (
	.Y(N18),
	.D(n8),
	.C(n9),
	.B(n10),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U26 (
	.Y(n29),
	.S0(\RX_IN_reg[0] ),
	.B(n16),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U27 (
	.Y(n12),
	.B(n16),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   MXI2X1M U28 (
	.Y(n28),
	.S0(N25),
	.B(n19),
	.A(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U29 (
	.Y(n19),
	.B0(n20),
	.A1N(\RX_IN_reg[0] ),
	.A0(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X1M U30 (
	.Y(n18),
	.C(n17),
	.B(n16),
	.A(\RX_IN_reg[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKINVX1M U31 (
	.Y(n16),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X1M U32 (
	.Y(n20),
	.B0(n22),
	.A1(n21),
	.A0(RX_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKMX2X2M U33 (
	.Y(n27),
	.S0(n22),
	.B(n23),
	.A(sample_bit_samp), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U34 (
	.Y(n22),
	.B0(n17),
	.A1N(N18),
	.A0(data_samp_en), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U35 (
	.Y(n17),
	.B(n21),
	.A(data_samp_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X1M U36 (
	.Y(n21),
	.C(n24),
	.B(edge_cnt[1]),
	.A(edge_cnt[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR3X1M U37 (
	.Y(n24),
	.C(edge_cnt[3]),
	.B(edge_cnt[4]),
	.A(edge_cnt[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U38 (
	.Y(n23),
	.B(data_samp_en),
	.AN(N25), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module edge_bit_counter_RX_test_1 (
	CLK_EDGE, 
	RST_EDGE, 
	enable_edge, 
	prescale_edge, 
	bit_cnt_edge, 
	edge_cnt_edge, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK_EDGE;
   input RST_EDGE;
   input enable_edge;
   input [5:0] prescale_edge;
   output [5:0] bit_cnt_edge;
   output [5:0] edge_cnt_edge;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N7;
   wire N8;
   wire N9;
   wire N10;
   wire N11;
   wire N12;
   wire N13;
   wire N15;
   wire N16;
   wire N17;
   wire N18;
   wire N19;
   wire N20;
   wire N28;
   wire N31;
   wire N32;
   wire N33;
   wire N34;
   wire N35;
   wire N42;
   wire N43;
   wire N44;
   wire N45;
   wire N46;
   wire N47;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire \add_32/carry[5] ;
   wire \add_32/carry[4] ;
   wire \add_32/carry[3] ;
   wire \add_32/carry[2] ;
   wire \add_16/carry[5] ;
   wire \add_16/carry[4] ;
   wire \add_16/carry[3] ;
   wire \add_16/carry[2] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;

   // Module instantiations
   SDFFRQX2M \bit_cnt_edge_reg[5]  (
	.SI(bit_cnt_edge[4]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(bit_cnt_edge[5]),
	.D(n26),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_cnt_edge_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(bit_cnt_edge[0]),
	.D(n25),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_cnt_edge_reg[3]  (
	.SI(bit_cnt_edge[2]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(bit_cnt_edge[3]),
	.D(n22),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_cnt_edge_reg[4]  (
	.SI(bit_cnt_edge[3]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(bit_cnt_edge[4]),
	.D(n21),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_cnt_edge_reg[1]  (
	.SI(N15),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(bit_cnt_edge[1]),
	.D(n24),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \bit_cnt_edge_reg[2]  (
	.SI(bit_cnt_edge[1]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(bit_cnt_edge[2]),
	.D(n23),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_edge_reg[5]  (
	.SI(edge_cnt_edge[4]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(edge_cnt_edge[5]),
	.D(N47),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_edge_reg[4]  (
	.SI(edge_cnt_edge[3]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(edge_cnt_edge[4]),
	.D(N46),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_edge_reg[3]  (
	.SI(edge_cnt_edge[2]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(edge_cnt_edge[3]),
	.D(N45),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_edge_reg[2]  (
	.SI(n35),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(edge_cnt_edge[2]),
	.D(N44),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_edge_reg[1]  (
	.SI(edge_cnt_edge[0]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(edge_cnt_edge[1]),
	.D(N43),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \edge_cnt_edge_reg[0]  (
	.SI(bit_cnt_edge[5]),
	.SE(test_se),
	.RN(RST_EDGE),
	.Q(edge_cnt_edge[0]),
	.D(N42),
	.CK(CLK_EDGE), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U7 (
	.Y(n20),
	.B(enable_edge),
	.A(N28), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U8 (
	.Y(n18),
	.B(N28),
	.A(enable_edge), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U17 (
	.Y(n19),
	.B(n18),
	.AN(enable_edge), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U18 (
	.Y(N43),
	.B(n20),
	.AN(N31), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U19 (
	.Y(N44),
	.B(n20),
	.AN(N32), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U20 (
	.Y(N45),
	.B(n20),
	.AN(N33), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U21 (
	.Y(N46),
	.B(n20),
	.AN(N34), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U22 (
	.Y(N42),
	.B(n20),
	.A(edge_cnt_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U23 (
	.Y(N47),
	.C(N28),
	.B(enable_edge),
	.A(N35), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U24 (
	.Y(n21),
	.B1(n19),
	.B0(N19),
	.A1(n18),
	.A0(bit_cnt_edge[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U25 (
	.Y(n22),
	.B1(n19),
	.B0(N18),
	.A1(n18),
	.A0(bit_cnt_edge[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U26 (
	.Y(n23),
	.B1(n19),
	.B0(N17),
	.A1(n18),
	.A0(bit_cnt_edge[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U27 (
	.Y(n24),
	.B1(n19),
	.B0(N16),
	.A1(n18),
	.A0(bit_cnt_edge[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U28 (
	.Y(n25),
	.B1(n19),
	.B0(N15),
	.A1(n18),
	.A0(bit_cnt_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(N15),
	.A(bit_cnt_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U30 (
	.Y(n26),
	.B1(n19),
	.B0(N20),
	.A1(n18),
	.A0(bit_cnt_edge[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U31 (
	.Y(N7),
	.A(prescale_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U32 (
	.Y(n35),
	.A(edge_cnt_edge[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U33 (
	.S(N17),
	.CO(\add_16/carry[3] ),
	.B(\add_16/carry[2] ),
	.A(bit_cnt_edge[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U34 (
	.S(N16),
	.CO(\add_16/carry[2] ),
	.B(bit_cnt_edge[0]),
	.A(bit_cnt_edge[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U35 (
	.S(N31),
	.CO(\add_32/carry[2] ),
	.B(edge_cnt_edge[0]),
	.A(edge_cnt_edge[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U36 (
	.S(N18),
	.CO(\add_16/carry[4] ),
	.B(\add_16/carry[3] ),
	.A(bit_cnt_edge[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U37 (
	.S(N32),
	.CO(\add_32/carry[3] ),
	.B(\add_32/carry[2] ),
	.A(edge_cnt_edge[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U38 (
	.S(N33),
	.CO(\add_32/carry[4] ),
	.B(\add_32/carry[3] ),
	.A(edge_cnt_edge[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U39 (
	.S(N19),
	.CO(\add_16/carry[5] ),
	.B(\add_16/carry[4] ),
	.A(bit_cnt_edge[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   ADDHX1M U40 (
	.S(N34),
	.CO(\add_32/carry[5] ),
	.B(\add_32/carry[4] ),
	.A(edge_cnt_edge[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U41 (
	.Y(n1),
	.B(N7),
	.AN(prescale_edge[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U42 (
	.Y(N8),
	.B0(n1),
	.A1N(prescale_edge[1]),
	.A0N(prescale_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U43 (
	.Y(n2),
	.B(prescale_edge[2]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U44 (
	.Y(N9),
	.B0(n2),
	.A1N(prescale_edge[2]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U45 (
	.Y(n3),
	.B(prescale_edge[3]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U46 (
	.Y(N10),
	.B0(n3),
	.A1N(prescale_edge[3]),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U47 (
	.Y(n4),
	.B(prescale_edge[4]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U48 (
	.Y(N11),
	.B0(n4),
	.A1N(prescale_edge[4]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U49 (
	.Y(N13),
	.B(prescale_edge[5]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U50 (
	.Y(N12),
	.B0(N13),
	.A1(prescale_edge[5]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U51 (
	.Y(N20),
	.B(bit_cnt_edge[5]),
	.A(\add_16/carry[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U52 (
	.Y(N35),
	.B(edge_cnt_edge[5]),
	.A(\add_32/carry[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U53 (
	.Y(n34),
	.B(edge_cnt_edge[3]),
	.A(N10), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U54 (
	.Y(n33),
	.B(edge_cnt_edge[2]),
	.A(N9), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U55 (
	.Y(n32),
	.B(edge_cnt_edge[4]),
	.A(N11), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U56 (
	.Y(n5),
	.B(edge_cnt_edge[0]),
	.A(prescale_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U57 (
	.Y(n30),
	.B1(n5),
	.B0(N8),
	.A1(n35),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKNAND2X2M U58 (
	.Y(n27),
	.B(prescale_edge[0]),
	.A(edge_cnt_edge[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U59 (
	.Y(n29),
	.B1(N8),
	.B0(n27),
	.A1(n35),
	.A0(n27), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U60 (
	.Y(n28),
	.B(edge_cnt_edge[5]),
	.A(N12), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4BX1M U61 (
	.Y(n31),
	.D(N13),
	.C(n28),
	.B(n29),
	.AN(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X1M U62 (
	.Y(N28),
	.D(n31),
	.C(n32),
	.B(n33),
	.A(n34), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FSM_RX_test_1 (
	CLK_FSM, 
	RST_FSM, 
	RX_IN, 
	bit_cnt_FSM, 
	edge_cnt_FSM, 
	PAR_EN_FSM, 
	par_err_FSM, 
	strt_glitch_FSM, 
	stp_err_FSM, 
	prescale_FSM, 
	par_chk_en_FSM, 
	strt_chk_en_FSM, 
	stp_chk_en_FSM, 
	enable_FSM, 
	data_samp_en_FSM, 
	data_valid_FSM, 
	deser_en_FSM, 
	test_si, 
	test_so, 
	test_se, 
	VDD, 
	VSS);
   input CLK_FSM;
   input RST_FSM;
   input RX_IN;
   input [5:0] bit_cnt_FSM;
   input [5:0] edge_cnt_FSM;
   input PAR_EN_FSM;
   input par_err_FSM;
   input strt_glitch_FSM;
   input stp_err_FSM;
   input [5:0] prescale_FSM;
   output par_chk_en_FSM;
   output strt_chk_en_FSM;
   output stp_chk_en_FSM;
   output enable_FSM;
   output data_samp_en_FSM;
   output data_valid_FSM;
   output deser_en_FSM;
   input test_si;
   output test_so;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire par_err_reg;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire \r107/EQ ;
   wire \r107/B[0] ;
   wire \r107/B[1] ;
   wire \r107/B[2] ;
   wire \r107/B[3] ;
   wire \r107/B[4] ;
   wire \r107/B[5] ;
   wire \r107/B[9] ;
   wire n1;
   wire n2;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n18;
   wire n19;
   wire n20;
   wire [2:0] cs;
   wire [2:0] ns;

   assign test_so = par_err_reg ;

   // Module instantiations
   SDFFRQX2M data_valid_FSM_reg (
	.SI(n19),
	.SE(test_se),
	.RN(RST_FSM),
	.Q(data_valid_FSM),
	.D(n60),
	.CK(CLK_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M par_err_reg_reg (
	.SI(data_valid_FSM),
	.SE(test_se),
	.RN(RST_FSM),
	.Q(par_err_reg),
	.D(n61),
	.CK(CLK_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cs_reg[2]  (
	.SI(n18),
	.SE(test_se),
	.RN(RST_FSM),
	.Q(cs[2]),
	.D(ns[2]),
	.CK(CLK_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cs_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_FSM),
	.Q(cs[0]),
	.D(ns[0]),
	.CK(CLK_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cs_reg[1]  (
	.SI(cs[0]),
	.SE(test_se),
	.RN(RST_FSM),
	.Q(cs[1]),
	.D(ns[1]),
	.CK(CLK_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n16),
	.A(n49), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U9 (
	.Y(n20),
	.A(\r107/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U10 (
	.Y(par_chk_en_FSM),
	.B(n44),
	.AN(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U11 (
	.Y(deser_en_FSM),
	.B(n54),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U12 (
	.Y(stp_chk_en_FSM),
	.C(n19),
	.B(n20),
	.A(n44), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U13 (
	.Y(n49),
	.B(n55),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U14 (
	.Y(data_samp_en_FSM),
	.B0(n44),
	.A1N(n59),
	.A0N(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U15 (
	.Y(n59),
	.B(n15),
	.A(RX_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U16 (
	.Y(n48),
	.B(cs[2]),
	.A(n20), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U17 (
	.Y(n50),
	.B0(n44),
	.A1(cs[2]),
	.A0(\r107/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U18 (
	.Y(enable_FSM),
	.B1(n58),
	.B0(cs[2]),
	.A1(n44),
	.A0(\r107/EQ ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U19 (
	.Y(n58),
	.B(n59),
	.A(cs[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BXLM U20 (
	.Y(n46),
	.D(n53),
	.C(bit_cnt_FSM[3]),
	.B(\r107/EQ ),
	.AN(bit_cnt_FSM[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U21 (
	.Y(n53),
	.D(bit_cnt_FSM[1]),
	.C(bit_cnt_FSM[2]),
	.B(bit_cnt_FSM[4]),
	.A(bit_cnt_FSM[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31XLM U22 (
	.Y(ns[2]),
	.B0(n45),
	.A2(n44),
	.A1(\r107/EQ ),
	.A0(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U23 (
	.Y(n45),
	.B0(par_chk_en_FSM),
	.A1N(n46),
	.A0(n47), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U24 (
	.Y(n47),
	.B(n16),
	.A(PAR_EN_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U25 (
	.Y(ns[1]),
	.C0(n16),
	.B0(n14),
	.A1(n43),
	.A0(strt_glitch_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U26 (
	.Y(n14),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X1M U27 (
	.Y(n55),
	.B(\r107/EQ ),
	.A(strt_glitch_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U28 (
	.Y(n61),
	.B1(n44),
	.B0(n57),
	.A1N(par_err_reg),
	.A0N(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U29 (
	.Y(n57),
	.B0(n44),
	.A1(n48),
	.A0(par_err_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B1X2M U30 (
	.Y(ns[0]),
	.B0(n51),
	.A1N(stp_chk_en_FSM),
	.A0(RX_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI32X1M U31 (
	.Y(n51),
	.B1(n46),
	.B0(n49),
	.A2(n52),
	.A1(n19),
	.A0(n18), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U32 (
	.Y(n52),
	.B1(n15),
	.B0(n55),
	.A1(RX_IN),
	.A0(cs[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U33 (
	.Y(n43),
	.C(cs[0]),
	.B(n18),
	.A(n48), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U34 (
	.Y(\r107/B[0] ),
	.A(prescale_FSM[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U35 (
	.Y(n60),
	.B0(n56),
	.A1(n50),
	.A0(data_valid_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U36 (
	.Y(n56),
	.D(n44),
	.C(n50),
	.B(par_err_reg),
	.A(stp_err_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U37 (
	.Y(strt_chk_en_FSM),
	.A(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U38 (
	.Y(n44),
	.B(n15),
	.A(cs[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U39 (
	.Y(n15),
	.A(cs[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U40 (
	.Y(n19),
	.A(cs[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U41 (
	.Y(n54),
	.C(cs[1]),
	.B(n19),
	.A(cs[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U42 (
	.Y(n18),
	.A(cs[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2BX1M U43 (
	.Y(n1),
	.B(\r107/B[0] ),
	.AN(prescale_FSM[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U44 (
	.Y(\r107/B[1] ),
	.B0(n1),
	.A1N(prescale_FSM[1]),
	.A0N(prescale_FSM[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U45 (
	.Y(n2),
	.B(prescale_FSM[2]),
	.A(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U46 (
	.Y(\r107/B[2] ),
	.B0(n2),
	.A1N(prescale_FSM[2]),
	.A0N(n1), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U47 (
	.Y(n3),
	.B(prescale_FSM[3]),
	.A(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U48 (
	.Y(\r107/B[3] ),
	.B0(n3),
	.A1N(prescale_FSM[3]),
	.A0N(n2), 
	.VDD(VDD), 
	.VSS(VSS));
   OR2X1M U49 (
	.Y(n4),
	.B(prescale_FSM[4]),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X1M U50 (
	.Y(\r107/B[4] ),
	.B0(n4),
	.A1N(prescale_FSM[4]),
	.A0N(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X1M U51 (
	.Y(\r107/B[9] ),
	.B(prescale_FSM[5]),
	.A(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U52 (
	.Y(\r107/B[5] ),
	.B0(\r107/B[9] ),
	.A1(prescale_FSM[5]),
	.A0(n4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U53 (
	.Y(n5),
	.B(edge_cnt_FSM[0]),
	.AN(\r107/B[0] ), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U54 (
	.Y(n9),
	.B1(n5),
	.B0(\r107/B[1] ),
	.A1N(edge_cnt_FSM[1]),
	.A0(n5), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X1M U55 (
	.Y(n8),
	.B(edge_cnt_FSM[5]),
	.A(\r107/B[5] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX1M U56 (
	.Y(n6),
	.B(\r107/B[0] ),
	.AN(edge_cnt_FSM[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U57 (
	.Y(n7),
	.B1(n6),
	.B0(edge_cnt_FSM[1]),
	.A1N(\r107/B[1] ),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U58 (
	.Y(n13),
	.D(n7),
	.C(n8),
	.B(n9),
	.AN(\r107/B[9] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U59 (
	.Y(n12),
	.B(edge_cnt_FSM[4]),
	.A(\r107/B[4] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U60 (
	.Y(n11),
	.B(edge_cnt_FSM[2]),
	.A(\r107/B[2] ), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U61 (
	.Y(n10),
	.B(edge_cnt_FSM[3]),
	.A(\r107/B[3] ), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U62 (
	.Y(\r107/EQ ),
	.D(n10),
	.C(n11),
	.B(n12),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module TOP_TX_DATA_LENGTH8_test_1 (
	RST, 
	CLK, 
	P_DATA, 
	PAR_TYP, 
	PAR_EN, 
	DATA_VALID, 
	TX_OUT, 
	BUSY, 
	test_si2, 
	test_si1, 
	test_so1, 
	test_se, 
	FE_OFN4_RST_SYNC_2_mux, 
	TX_CLK_M__L3_N2, 
	TX_CLK_M__L3_N3, 
	VDD, 
	VSS);
   input RST;
   input CLK;
   input [7:0] P_DATA;
   input PAR_TYP;
   input PAR_EN;
   input DATA_VALID;
   output TX_OUT;
   output BUSY;
   input test_si2;
   input test_si1;
   output test_so1;
   input test_se;
   input FE_OFN4_RST_SYNC_2_mux;
   input TX_CLK_M__L3_N2;
   input TX_CLK_M__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire ser_data;
   wire par_bit;
   wire ser_en;
   wire ser_done;
   wire n2;
   wire n3;
   wire [1:0] mux_sel;

   // Module instantiations
   MUX4x1_test_1 mux (
	.CLK_mux(TX_CLK_M__L3_N2),
	.RST_mux(RST),
	.start_bit_mux(1'b0),
	.stop_bit_mux(1'b1),
	.ser_data_mux(ser_data),
	.parity_bit_mux(par_bit),
	.mux_sel_mux({ mux_sel[1],
		mux_sel[0] }),
	.TX_OUT_mux(TX_OUT),
	.test_si(test_si2),
	.test_se(test_se), 
	.VDD(VDD), 
	.VSS(VSS));
   parity_calc_DATA_LENGTH8_test_1 PAR (
	.CLK(CLK),
	.RST(RST),
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.PAR_TYP(PAR_TYP),
	.Data_Valid(DATA_VALID),
	.PAR_EN(PAR_EN),
	.busy(BUSY),
	.par_bit(par_bit),
	.test_si(n3),
	.test_so(n2),
	.test_se(test_se),
	.FE_OFN4_RST_SYNC_2_mux(FE_OFN4_RST_SYNC_2_mux),
	.TX_CLK_M__L3_N2(TX_CLK_M__L3_N2),
	.TX_CLK_M__L3_N3(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SERIALIZER_DATA_LENGTH8_test_1 SER (
	.P_DATA({ P_DATA[7],
		P_DATA[6],
		P_DATA[5],
		P_DATA[4],
		P_DATA[3],
		P_DATA[2],
		P_DATA[1],
		P_DATA[0] }),
	.ser_en(ser_en),
	.CLK(TX_CLK_M__L3_N2),
	.RST(RST),
	.Data_Valid(DATA_VALID),
	.busy(BUSY),
	.ser_done(ser_done),
	.ser_data(ser_data),
	.test_si(n2),
	.test_so(test_so1),
	.test_se(test_se),
	.FE_OFN4_RST_SYNC_2_mux(FE_OFN4_RST_SYNC_2_mux),
	.TX_CLK_M__L3_N3(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   FSM_TX_test_1 FSM1 (
	.DATA_VALID_FSM(DATA_VALID),
	.RST_FSM(RST),
	.CLK_FSM(CLK),
	.SER_DONE_FSM(ser_done),
	.PAR_EN_FSM(PAR_EN),
	.SER_EN_FSM(ser_en),
	.BUSY_FSM(BUSY),
	.MUX_SEL_FSM({ mux_sel[1],
		mux_sel[0] }),
	.test_si(test_si1),
	.test_so(n3),
	.test_se(test_se),
	.FE_OFN4_RST_SYNC_2_mux(FE_OFN4_RST_SYNC_2_mux),
	.TX_CLK_M__L3_N2(TX_CLK_M__L3_N2),
	.TX_CLK_M__L3_N3(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module MUX4x1_test_1 (
	CLK_mux, 
	RST_mux, 
	start_bit_mux, 
	stop_bit_mux, 
	ser_data_mux, 
	parity_bit_mux, 
	mux_sel_mux, 
	TX_OUT_mux, 
	test_si, 
	test_se, 
	VDD, 
	VSS);
   input CLK_mux;
   input RST_mux;
   input start_bit_mux;
   input stop_bit_mux;
   input ser_data_mux;
   input parity_bit_mux;
   input [1:0] mux_sel_mux;
   output TX_OUT_mux;
   input test_si;
   input test_se;
   inout VDD;
   inout VSS;

   // Internal wires
   wire HTIE_LTIEHI_NET;
   wire LTIE_LTIELO_NET;
   wire TX_OUT_mux_c;
   wire n3;
   wire n4;
   wire n2;

   // Module instantiations
   TIEHIM HTIE_LTIEHI (
	.Y(HTIE_LTIEHI_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   TIELOM LTIE_LTIELO (
	.Y(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M TX_OUT_mux_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_mux),
	.Q(TX_OUT_mux),
	.D(TX_OUT_mux_c),
	.CK(CLK_mux), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U4 (
	.Y(n2),
	.A(mux_sel_mux[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2B2X1M U5 (
	.Y(TX_OUT_mux_c),
	.B1(n4),
	.B0(mux_sel_mux[1]),
	.A1N(mux_sel_mux[1]),
	.A0(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U6 (
	.Y(n4),
	.B1(mux_sel_mux[0]),
	.B0(HTIE_LTIEHI_NET),
	.A1(n2),
	.A0(LTIE_LTIELO_NET), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U7 (
	.Y(n3),
	.B1(mux_sel_mux[0]),
	.B0(parity_bit_mux),
	.A1(n2),
	.A0(ser_data_mux), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module parity_calc_DATA_LENGTH8_test_1 (
	CLK, 
	RST, 
	P_DATA, 
	PAR_TYP, 
	Data_Valid, 
	PAR_EN, 
	busy, 
	par_bit, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN4_RST_SYNC_2_mux, 
	TX_CLK_M__L3_N2, 
	TX_CLK_M__L3_N3, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [7:0] P_DATA;
   input PAR_TYP;
   input Data_Valid;
   input PAR_EN;
   input busy;
   output par_bit;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN4_RST_SYNC_2_mux;
   input TX_CLK_M__L3_N2;
   input TX_CLK_M__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire n1;
   wire n3;
   wire n4;
   wire n5;
   wire n6;
   wire n7;
   wire n9;
   wire n11;
   wire n13;
   wire n15;
   wire n17;
   wire n19;
   wire n21;
   wire n23;
   wire n25;
   wire n2;
   wire [7:0] par_data;

   assign test_so = par_data[7] ;

   // Module instantiations
   SDFFRQX2M \par_data_reg[5]  (
	.SI(par_data[4]),
	.SE(test_se),
	.RN(RST),
	.Q(par_data[5]),
	.D(n21),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \par_data_reg[1]  (
	.SI(par_data[0]),
	.SE(test_se),
	.RN(RST),
	.Q(par_data[1]),
	.D(n13),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \par_data_reg[4]  (
	.SI(par_data[3]),
	.SE(test_se),
	.RN(RST),
	.Q(par_data[4]),
	.D(n19),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \par_data_reg[0]  (
	.SI(par_bit),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(par_data[0]),
	.D(n11),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \par_data_reg[2]  (
	.SI(par_data[1]),
	.SE(test_se),
	.RN(RST),
	.Q(par_data[2]),
	.D(n15),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M par_bit_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(par_bit),
	.D(n9),
	.CK(TX_CLK_M__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \par_data_reg[3]  (
	.SI(par_data[2]),
	.SE(test_se),
	.RN(RST),
	.Q(par_data[3]),
	.D(n17),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \par_data_reg[6]  (
	.SI(par_data[5]),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(par_data[6]),
	.D(n23),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \par_data_reg[7]  (
	.SI(par_data[6]),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(par_data[7]),
	.D(n25),
	.CK(TX_CLK_M__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U2 (
	.Y(n7),
	.B(busy),
	.AN(Data_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U3 (
	.Y(n11),
	.B1(n7),
	.B0(P_DATA[0]),
	.A1N(n7),
	.A0(par_data[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U4 (
	.Y(n13),
	.B1(n7),
	.B0(P_DATA[1]),
	.A1N(n7),
	.A0(par_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U5 (
	.Y(n15),
	.B1(n7),
	.B0(P_DATA[2]),
	.A1N(n7),
	.A0(par_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U6 (
	.Y(n17),
	.B1(n7),
	.B0(P_DATA[3]),
	.A1N(n7),
	.A0(par_data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U7 (
	.Y(n19),
	.B1(n7),
	.B0(P_DATA[4]),
	.A1N(n7),
	.A0(par_data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U8 (
	.Y(n21),
	.B1(n7),
	.B0(P_DATA[5]),
	.A1N(n7),
	.A0(par_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U9 (
	.Y(n23),
	.B1(n7),
	.B0(P_DATA[6]),
	.A1N(n7),
	.A0(par_data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO2B2X2M U10 (
	.Y(n25),
	.B1(n7),
	.B0(P_DATA[7]),
	.A1N(n7),
	.A0(par_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U11 (
	.Y(n5),
	.B(par_data[3]),
	.A(par_data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U12 (
	.Y(n3),
	.C(n6),
	.B(par_data[4]),
	.A(par_data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   CLKXOR2X2M U13 (
	.Y(n6),
	.B(par_data[6]),
	.A(par_data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U14 (
	.Y(n9),
	.B1(n2),
	.B0(n1),
	.A1N(n2),
	.A0N(par_bit), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n2),
	.A(PAR_EN), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U16 (
	.Y(n1),
	.C(n4),
	.B(PAR_TYP),
	.A(n3), 
	.VDD(VDD), 
	.VSS(VSS));
   XOR3XLM U17 (
	.Y(n4),
	.C(n5),
	.B(par_data[0]),
	.A(par_data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SERIALIZER_DATA_LENGTH8_test_1 (
	P_DATA, 
	ser_en, 
	CLK, 
	RST, 
	Data_Valid, 
	busy, 
	ser_done, 
	ser_data, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN4_RST_SYNC_2_mux, 
	TX_CLK_M__L3_N3, 
	VDD, 
	VSS);
   input [7:0] P_DATA;
   input ser_en;
   input CLK;
   input RST;
   input Data_Valid;
   input busy;
   output ser_done;
   output ser_data;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN4_RST_SYNC_2_mux;
   input TX_CLK_M__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire N24;
   wire N25;
   wire N26;
   wire N27;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n13;
   wire n14;
   wire n15;
   wire [7:1] data;
   wire [3:0] counter;

   assign test_so = data[7] ;

   // Module instantiations
   SDFFSQX2M \data_reg[6]  (
	.SN(RST),
	.SI(data[5]),
	.SE(test_se),
	.Q(data[6]),
	.D(n32),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \data_reg[5]  (
	.SN(FE_OFN4_RST_SYNC_2_mux),
	.SI(data[4]),
	.SE(test_se),
	.Q(data[5]),
	.D(n33),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \data_reg[4]  (
	.SN(FE_OFN4_RST_SYNC_2_mux),
	.SI(data[3]),
	.SE(test_se),
	.Q(data[4]),
	.D(n34),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \data_reg[3]  (
	.SN(FE_OFN4_RST_SYNC_2_mux),
	.SI(data[2]),
	.SE(test_se),
	.Q(data[3]),
	.D(n35),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \data_reg[2]  (
	.SN(FE_OFN4_RST_SYNC_2_mux),
	.SI(data[1]),
	.SE(test_se),
	.Q(data[2]),
	.D(n36),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \data_reg[1]  (
	.SN(FE_OFN4_RST_SYNC_2_mux),
	.SI(ser_data),
	.SE(test_se),
	.Q(data[1]),
	.D(n37),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \data_reg[0]  (
	.SN(FE_OFN4_RST_SYNC_2_mux),
	.SI(counter[3]),
	.SE(test_se),
	.Q(ser_data),
	.D(n30),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFSQX2M \data_reg[7]  (
	.SN(FE_OFN4_RST_SYNC_2_mux),
	.SI(data[6]),
	.SE(test_se),
	.Q(data[7]),
	.D(n31),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[3]  (
	.SI(n14),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(counter[3]),
	.D(N27),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[1]  (
	.SI(counter[0]),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(counter[1]),
	.D(N25),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[2]  (
	.SI(counter[1]),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(counter[2]),
	.D(N26),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \counter_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(counter[0]),
	.D(N24),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U15 (
	.Y(n18),
	.B(n19),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U16 (
	.Y(n16),
	.B(n18),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n13),
	.A(ser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U18 (
	.Y(n19),
	.B(busy),
	.AN(Data_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U19 (
	.Y(n30),
	.B0(n17),
	.A1N(n16),
	.A0N(ser_data), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U20 (
	.Y(n17),
	.B1(n19),
	.B0(P_DATA[0]),
	.A1(n18),
	.A0(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U21 (
	.Y(n37),
	.B0(n25),
	.A1N(n16),
	.A0N(data[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U22 (
	.Y(n25),
	.B1(n19),
	.B0(P_DATA[1]),
	.A1(n18),
	.A0(data[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U23 (
	.Y(n36),
	.B0(n24),
	.A1N(data[2]),
	.A0N(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U24 (
	.Y(n24),
	.B1(n19),
	.B0(P_DATA[2]),
	.A1(n18),
	.A0(data[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U25 (
	.Y(n35),
	.B0(n23),
	.A1N(data[3]),
	.A0N(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U26 (
	.Y(n23),
	.B1(n19),
	.B0(P_DATA[3]),
	.A1(n18),
	.A0(data[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U27 (
	.Y(n34),
	.B0(n22),
	.A1N(data[4]),
	.A0N(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U28 (
	.Y(n22),
	.B1(n19),
	.B0(P_DATA[4]),
	.A1(n18),
	.A0(data[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U29 (
	.Y(n33),
	.B0(n21),
	.A1N(data[5]),
	.A0N(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U30 (
	.Y(n21),
	.B1(n19),
	.B0(P_DATA[5]),
	.A1(n18),
	.A0(data[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U31 (
	.Y(n32),
	.B0(n20),
	.A1N(data[6]),
	.A0N(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U32 (
	.Y(n20),
	.B1(n19),
	.B0(P_DATA[6]),
	.A1(n18),
	.A0(data[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AO22X1M U33 (
	.Y(n31),
	.B1(n19),
	.B0(P_DATA[7]),
	.A1(data[7]),
	.A0(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U34 (
	.Y(N27),
	.B1(n15),
	.B0(n27),
	.A2(n26),
	.A1(counter[3]),
	.A0(n14), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U35 (
	.Y(n27),
	.B0(n28),
	.A1(counter[2]),
	.A0(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U36 (
	.Y(ser_done),
	.D(n15),
	.C(counter[0]),
	.B(counter[1]),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI2B1X1M U37 (
	.Y(n28),
	.B0(N24),
	.A1N(counter[1]),
	.A0(ser_en), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U38 (
	.Y(n26),
	.C(counter[1]),
	.B(ser_en),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U39 (
	.Y(N26),
	.B1(n26),
	.B0(counter[2]),
	.A1(n14),
	.A0(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U40 (
	.Y(N24),
	.B(counter[0]),
	.A(n13), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U41 (
	.Y(N25),
	.B(n13),
	.A(n29), 
	.VDD(VDD), 
	.VSS(VSS));
   XNOR2X2M U42 (
	.Y(n29),
	.B(counter[1]),
	.A(counter[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U43 (
	.Y(n15),
	.A(counter[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U44 (
	.Y(n14),
	.A(counter[2]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module FSM_TX_test_1 (
	DATA_VALID_FSM, 
	RST_FSM, 
	CLK_FSM, 
	SER_DONE_FSM, 
	PAR_EN_FSM, 
	SER_EN_FSM, 
	BUSY_FSM, 
	MUX_SEL_FSM, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN4_RST_SYNC_2_mux, 
	TX_CLK_M__L3_N2, 
	TX_CLK_M__L3_N3, 
	VDD, 
	VSS);
   input DATA_VALID_FSM;
   input RST_FSM;
   input CLK_FSM;
   input SER_DONE_FSM;
   input PAR_EN_FSM;
   output SER_EN_FSM;
   output BUSY_FSM;
   output [1:0] MUX_SEL_FSM;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN4_RST_SYNC_2_mux;
   input TX_CLK_M__L3_N2;
   input TX_CLK_M__L3_N3;
   inout VDD;
   inout VSS;

   // Internal wires
   wire BUSY_FSM_c;
   wire n11;
   wire n12;
   wire n13;
   wire n5;
   wire n6;
   wire n7;
   wire n8;
   wire n9;
   wire n10;
   wire [2:0] cs;
   wire [2:0] ns;

   assign test_so = n8 ;

   // Module instantiations
   SDFFRQX2M BUSY_FSM_reg (
	.SI(test_si),
	.SE(test_se),
	.RN(RST_FSM),
	.Q(BUSY_FSM),
	.D(BUSY_FSM_c),
	.CK(CLK_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cs_reg[0]  (
	.SI(BUSY_FSM),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(cs[0]),
	.D(ns[0]),
	.CK(TX_CLK_M__L3_N3), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cs_reg[2]  (
	.SI(cs[1]),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(cs[2]),
	.D(ns[2]),
	.CK(TX_CLK_M__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \cs_reg[1]  (
	.SI(n6),
	.SE(test_se),
	.RN(FE_OFN4_RST_SYNC_2_mux),
	.Q(cs[1]),
	.D(ns[1]),
	.CK(TX_CLK_M__L3_N2), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U7 (
	.Y(SER_EN_FSM),
	.B1(n11),
	.B0(SER_DONE_FSM),
	.A2(cs[1]),
	.A1(cs[2]),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U8 (
	.Y(n10),
	.A(DATA_VALID_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U9 (
	.Y(MUX_SEL_FSM[0]),
	.C(n13),
	.B(n8),
	.A(n12), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U10 (
	.Y(n13),
	.B1(n6),
	.B0(n10),
	.A1(n7),
	.A0(SER_DONE_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   AO21XLM U11 (
	.Y(BUSY_FSM_c),
	.B0(ns[1]),
	.A1(DATA_VALID_FSM),
	.A0(n8), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U12 (
	.Y(n5),
	.A(SER_EN_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U13 (
	.Y(n7),
	.A(n11), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI31X1M U14 (
	.Y(ns[0]),
	.B0(n5),
	.A2(cs[1]),
	.A1(cs[2]),
	.A0(n10), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U15 (
	.Y(MUX_SEL_FSM[1]),
	.B0(n5),
	.A1N(PAR_EN_FSM),
	.A0N(n7), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U16 (
	.Y(n11),
	.C(cs[1]),
	.B(n8),
	.A(cs[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U17 (
	.Y(n8),
	.A(cs[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n6),
	.A(cs[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI32X1M U19 (
	.Y(ns[2]),
	.B1(n12),
	.B0(cs[2]),
	.A2(n11),
	.A1(PAR_EN_FSM),
	.A0(n9), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n9),
	.A(SER_DONE_FSM), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U21 (
	.Y(ns[1]),
	.B0(cs[2]),
	.A1(n12),
	.A0(n6), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U22 (
	.Y(n12),
	.B(n6),
	.A(cs[1]), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_CTRL_test_1 (
	CLK, 
	RST, 
	ALU_OUT, 
	OUT_Valid, 
	CTRL_FULL_IN, 
	RdData, 
	RdData_Valid, 
	RX_P_DATA, 
	RX_D_VLD, 
	ALU_FUN, 
	ALU_EN, 
	CLK_EN, 
	Address, 
	WrEn, 
	RdEn, 
	WrData, 
	TX_P_DATA, 
	TX_D_VLD, 
	clk_div_en, 
	test_si, 
	test_so, 
	test_se, 
	FE_OFN0_RST_SYNC_1_mux, 
	CLK_R_M__L5_N4, 
	VDD, 
	VSS);
   input CLK;
   input RST;
   input [15:0] ALU_OUT;
   input OUT_Valid;
   input CTRL_FULL_IN;
   input [7:0] RdData;
   input RdData_Valid;
   input [7:0] RX_P_DATA;
   input RX_D_VLD;
   output [3:0] ALU_FUN;
   output ALU_EN;
   output CLK_EN;
   output [3:0] Address;
   output WrEn;
   output RdEn;
   output [7:0] WrData;
   output [7:0] TX_P_DATA;
   output TX_D_VLD;
   output clk_div_en;
   input test_si;
   output test_so;
   input test_se;
   input FE_OFN0_RST_SYNC_1_mux;
   input CLK_R_M__L5_N4;
   inout VDD;
   inout VSS;

   // Internal wires
   wire second_frame;
   wire second_frame_reg;
   wire n28;
   wire n29;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire n45;
   wire n46;
   wire n47;
   wire n48;
   wire n49;
   wire n50;
   wire n51;
   wire n52;
   wire n53;
   wire n54;
   wire n55;
   wire n56;
   wire n57;
   wire n58;
   wire n59;
   wire n60;
   wire n61;
   wire n62;
   wire n63;
   wire n64;
   wire n65;
   wire n66;
   wire n67;
   wire n68;
   wire n69;
   wire n70;
   wire n71;
   wire n72;
   wire n73;
   wire n74;
   wire n75;
   wire n76;
   wire n77;
   wire n78;
   wire n79;
   wire n80;
   wire n81;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n16;
   wire n17;
   wire n18;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n23;
   wire n24;
   wire n25;
   wire n26;
   wire n27;
   wire n82;
   wire [3:0] current_state;
   wire [3:0] next_state;

   assign clk_div_en = 1'b1 ;
   assign test_so = second_frame ;

   // Module instantiations
   SDFFRQX2M \Address_reg[2]  (
	.SI(Address[1]),
	.SE(test_se),
	.RN(RST),
	.Q(Address[2]),
	.D(n80),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Address_reg[3]  (
	.SI(Address[2]),
	.SE(test_se),
	.RN(RST),
	.Q(Address[3]),
	.D(n81),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \Address_reg[0]  (
	.SI(test_si),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(Address[0]),
	.D(n78),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX4M \Address_reg[1]  (
	.SI(Address[0]),
	.SE(test_se),
	.RN(RST),
	.Q(Address[1]),
	.D(n79),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M second_frame_reg_inst (
	.SI(n19),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(second_frame),
	.D(second_frame_reg),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[2]  (
	.SI(n22),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(current_state[2]),
	.D(next_state[2]),
	.CK(CLK), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[1]  (
	.SI(n16),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[1]),
	.D(next_state[1]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[0]  (
	.SI(Address[3]),
	.SE(test_se),
	.RN(RST),
	.Q(current_state[0]),
	.D(next_state[0]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   SDFFRQX2M \current_state_reg[3]  (
	.SI(n20),
	.SE(test_se),
	.RN(FE_OFN0_RST_SYNC_1_mux),
	.Q(current_state[3]),
	.D(next_state[3]),
	.CK(CLK_R_M__L5_N4), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U12 (
	.Y(ALU_FUN[2]),
	.B(n62),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U13 (
	.Y(ALU_EN),
	.B1(n55),
	.B0(OUT_Valid),
	.A1(n54),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U14 (
	.Y(WrData[0]),
	.B(n23),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U15 (
	.Y(n14),
	.A(WrEn), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U16 (
	.Y(n21),
	.A(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U17 (
	.Y(n59),
	.B(n31),
	.A(n15), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U18 (
	.Y(n23),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U19 (
	.Y(n15),
	.A(n61), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U20 (
	.Y(n12),
	.A(n55), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U21 (
	.Y(ALU_FUN[0]),
	.B(n54),
	.A(n23), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U22 (
	.Y(n64),
	.C0(n31),
	.B0(n18),
	.A1(n46),
	.A0(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U23 (
	.Y(n18),
	.A(n66), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U24 (
	.Y(n31),
	.C(n19),
	.B(current_state[2]),
	.A(n17), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U25 (
	.Y(WrEn),
	.B(n64),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U26 (
	.Y(n68),
	.B(n56),
	.A(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U27 (
	.Y(n46),
	.B(current_state[2]),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U28 (
	.Y(n17),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U29 (
	.Y(n11),
	.A(CTRL_FULL_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   OR3X2M U30 (
	.Y(TX_D_VLD),
	.C(n68),
	.B(second_frame_reg),
	.A(n69), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U31 (
	.Y(WrData[1]),
	.B(n58),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U32 (
	.Y(WrData[2]),
	.B(n62),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2XLM U33 (
	.Y(WrData[3]),
	.B(n63),
	.A(n64), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U34 (
	.Y(WrData[4]),
	.B(n14),
	.A(n26), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U35 (
	.Y(WrData[6]),
	.B(n14),
	.A(n25), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U36 (
	.Y(n39),
	.B0(n12),
	.A1(n13),
	.A0(n50), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U37 (
	.Y(next_state[0]),
	.D(n53),
	.C(n52),
	.B(n43),
	.A(n51), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U38 (
	.Y(n52),
	.C(n57),
	.B(n20),
	.A(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4BX1M U39 (
	.Y(n51),
	.D(n26),
	.C(n82),
	.B(n49),
	.AN(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   OA21X2M U40 (
	.Y(n53),
	.B0(n39),
	.A1(n24),
	.A0(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U41 (
	.Y(n61),
	.B(n34),
	.AN(n43), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U42 (
	.Y(n54),
	.C(n65),
	.B(n19),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U43 (
	.Y(n40),
	.B(n24),
	.A(n82), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U44 (
	.Y(n55),
	.C(current_state[2]),
	.B(n22),
	.A(n57), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U45 (
	.Y(n43),
	.C(n57),
	.B(n20),
	.A(n22), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U46 (
	.Y(n20),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U47 (
	.Y(n13),
	.A(n56), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U48 (
	.Y(ALU_FUN[1]),
	.B(n54),
	.A(n58), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U49 (
	.Y(ALU_FUN[3]),
	.B(n63),
	.A(n54), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U50 (
	.Y(n57),
	.B(current_state[3]),
	.A(n16), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2X2M U51 (
	.Y(n65),
	.B(current_state[0]),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U52 (
	.Y(n69),
	.C(RdData_Valid),
	.B(n11),
	.A(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U53 (
	.Y(n19),
	.A(current_state[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U55 (
	.Y(n66),
	.C(current_state[3]),
	.B(current_state[2]),
	.A(n65), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U56 (
	.Y(n50),
	.B(n11),
	.A(second_frame), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U57 (
	.Y(n22),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U58 (
	.Y(n16),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U59 (
	.Y(second_frame_reg),
	.C(n56),
	.B(second_frame),
	.A(CTRL_FULL_IN), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U60 (
	.Y(n77),
	.C(n21),
	.B(current_state[0]),
	.A(n19), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U61 (
	.Y(n36),
	.C(n17),
	.B(current_state[3]),
	.A(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR2BX2M U62 (
	.Y(RdEn),
	.B(RdData_Valid),
	.AN(n77), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U63 (
	.Y(TX_P_DATA[0]),
	.B0(n76),
	.A1N(second_frame_reg),
	.A0N(ALU_OUT[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U64 (
	.Y(n76),
	.B1(n69),
	.B0(RdData[0]),
	.A1(n68),
	.A0(ALU_OUT[8]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U65 (
	.Y(TX_P_DATA[1]),
	.B0(n75),
	.A1N(second_frame_reg),
	.A0N(ALU_OUT[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U66 (
	.Y(n75),
	.B1(n69),
	.B0(RdData[1]),
	.A1(n68),
	.A0(ALU_OUT[9]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U67 (
	.Y(TX_P_DATA[2]),
	.B0(n74),
	.A1N(second_frame_reg),
	.A0N(ALU_OUT[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U68 (
	.Y(n74),
	.B1(n69),
	.B0(RdData[2]),
	.A1(n68),
	.A0(ALU_OUT[10]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U69 (
	.Y(TX_P_DATA[3]),
	.B0(n73),
	.A1N(second_frame_reg),
	.A0N(ALU_OUT[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U70 (
	.Y(n73),
	.B1(n69),
	.B0(RdData[3]),
	.A1(n68),
	.A0(ALU_OUT[11]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U71 (
	.Y(TX_P_DATA[4]),
	.B0(n72),
	.A1N(second_frame_reg),
	.A0N(ALU_OUT[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U72 (
	.Y(n72),
	.B1(n69),
	.B0(RdData[4]),
	.A1(n68),
	.A0(ALU_OUT[12]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U73 (
	.Y(TX_P_DATA[5]),
	.B0(n71),
	.A1N(second_frame_reg),
	.A0N(ALU_OUT[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U74 (
	.Y(n71),
	.B1(n69),
	.B0(RdData[5]),
	.A1(n68),
	.A0(ALU_OUT[13]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U75 (
	.Y(TX_P_DATA[6]),
	.B0(n70),
	.A1N(second_frame_reg),
	.A0N(ALU_OUT[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U76 (
	.Y(n70),
	.B1(n69),
	.B0(RdData[6]),
	.A1(n68),
	.A0(ALU_OUT[14]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U77 (
	.Y(TX_P_DATA[7]),
	.B0(n67),
	.A1N(second_frame_reg),
	.A0N(ALU_OUT[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U78 (
	.Y(n67),
	.B1(n69),
	.B0(RdData[7]),
	.A1(n68),
	.A0(ALU_OUT[15]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U79 (
	.Y(n24),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U80 (
	.Y(next_state[2]),
	.C0(n39),
	.B0(n38),
	.A1(n17),
	.A0(n37), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U81 (
	.Y(n37),
	.B0(current_state[2]),
	.A1(current_state[3]),
	.A0(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND4X2M U82 (
	.Y(n38),
	.D(n42),
	.C(RX_P_DATA[4]),
	.B(n41),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U83 (
	.Y(n42),
	.D(n25),
	.C(n27),
	.B(RX_P_DATA[1]),
	.A(RX_P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI211X2M U84 (
	.Y(next_state[1]),
	.C0(n45),
	.B0(n44),
	.A1(n43),
	.A0(n24), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI211X2M U85 (
	.Y(n45),
	.C0(n48),
	.B0(n34),
	.A1(n47),
	.A0(n46), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U86 (
	.Y(n44),
	.B1(n50),
	.B0(n13),
	.A1(n12),
	.A0(OUT_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U87 (
	.Y(n47),
	.B1(RX_D_VLD),
	.B0(current_state[3]),
	.A1(RdData_Valid),
	.A0(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND3X2M U88 (
	.Y(n56),
	.C(current_state[2]),
	.B(n57),
	.A(current_state[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U89 (
	.Y(WrData[5]),
	.B(WrEn),
	.A(RX_P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND2X2M U90 (
	.Y(WrData[7]),
	.B(WrEn),
	.A(RX_P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND3X2M U91 (
	.Y(n41),
	.C(n36),
	.B(RX_P_DATA[3]),
	.A(RX_P_DATA[7]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U92 (
	.Y(n49),
	.D(n25),
	.C(n27),
	.B(n41),
	.A(RX_P_DATA[5]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U93 (
	.Y(n48),
	.D(RX_P_DATA[1]),
	.C(n49),
	.B(RX_P_DATA[4]),
	.A(n40), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR3X2M U94 (
	.Y(n34),
	.C(n21),
	.B(current_state[3]),
	.A(current_state[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   NOR4X1M U95 (
	.Y(n33),
	.D(RX_P_DATA[4]),
	.C(RX_P_DATA[5]),
	.B(RX_P_DATA[1]),
	.A(n35), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U96 (
	.Y(n35),
	.B(n82),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U97 (
	.Y(n63),
	.B(RX_P_DATA[3]),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U98 (
	.Y(n62),
	.B(RX_P_DATA[2]),
	.A(RX_D_VLD), 
	.VDD(VDD), 
	.VSS(VSS));
   NAND2X2M U99 (
	.Y(n58),
	.B(RX_D_VLD),
	.A(RX_P_DATA[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U100 (
	.Y(n79),
	.B1(n58),
	.B0(n61),
	.A1N(n59),
	.A0N(Address[1]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U101 (
	.Y(n80),
	.B1(n62),
	.B0(n61),
	.A1N(n59),
	.A0N(Address[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB2X1M U102 (
	.Y(n81),
	.B1(n63),
	.B0(n61),
	.A1N(n59),
	.A0N(Address[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI21X2M U103 (
	.Y(next_state[3]),
	.B0(n29),
	.A1(n24),
	.A0(n28), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI31X2M U104 (
	.Y(n29),
	.B0(n31),
	.A2(current_state[3]),
	.A1(n16),
	.A0(n30), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI21X2M U105 (
	.Y(n28),
	.B0(n34),
	.A1(n33),
	.A0(n32), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI22X1M U106 (
	.Y(n30),
	.B1(RX_D_VLD),
	.B0(current_state[1]),
	.A1(RdData_Valid),
	.A0(current_state[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U107 (
	.Y(n27),
	.A(RX_P_DATA[2]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U108 (
	.Y(n25),
	.A(RX_P_DATA[6]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U109 (
	.Y(n26),
	.A(RX_P_DATA[4]), 
	.VDD(VDD), 
	.VSS(VSS));
   AND4X2M U110 (
	.Y(n32),
	.D(n36),
	.C(RX_P_DATA[7]),
	.B(RX_P_DATA[6]),
	.A(RX_P_DATA[3]), 
	.VDD(VDD), 
	.VSS(VSS));
   INVX2M U111 (
	.Y(n82),
	.A(RX_P_DATA[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI2BB1X2M U112 (
	.Y(n78),
	.B0(n60),
	.A1N(n59),
	.A0N(Address[0]), 
	.VDD(VDD), 
	.VSS(VSS));
   AOI22X1M U113 (
	.Y(n60),
	.B1(n15),
	.B0(n40),
	.A1(RX_D_VLD),
	.A0(n31), 
	.VDD(VDD), 
	.VSS(VSS));
   OAI221X1M U114 (
	.Y(CLK_EN),
	.C0(n54),
	.B1(n66),
	.B0(n24),
	.A1(n55),
	.A0(OUT_Valid), 
	.VDD(VDD), 
	.VSS(VSS));
endmodule

module SYS_TOP (
	scan_clk, 
	scan_rst, 
	test_mode, 
	SE, 
	SI, 
	SO, 
	RST_N, 
	UART_CLK, 
	REF_CLK, 
	UART_RX_IN, 
	UART_TX_O, 
	parity_error, 
	framing_error, 
	VDD, 
	VSS);
   input scan_clk;
   input scan_rst;
   input test_mode;
   input SE;
   input [4:0] SI;
   output [4:0] SO;
   input RST_N;
   input UART_CLK;
   input REF_CLK;
   input UART_RX_IN;
   output UART_TX_O;
   output parity_error;
   output framing_error;
   inout VDD;
   inout VSS;

   // Internal wires
   wire REF_CLK__L2_N0;
   wire REF_CLK__L1_N0;
   wire UART_CLK__L2_N0;
   wire UART_CLK__L1_N0;
   wire scan_clk__L9_N0;
   wire scan_clk__L8_N1;
   wire scan_clk__L8_N0;
   wire scan_clk__L7_N0;
   wire scan_clk__L6_N0;
   wire scan_clk__L5_N0;
   wire scan_clk__L4_N0;
   wire scan_clk__L3_N0;
   wire scan_clk__L2_N1;
   wire scan_clk__L2_N0;
   wire scan_clk__L1_N0;
   wire CLK_R_M__L5_N7;
   wire CLK_R_M__L5_N6;
   wire CLK_R_M__L5_N5;
   wire CLK_R_M__L5_N4;
   wire CLK_R_M__L5_N3;
   wire CLK_R_M__L5_N2;
   wire CLK_R_M__L5_N1;
   wire CLK_R_M__L5_N0;
   wire CLK_R_M__L4_N3;
   wire CLK_R_M__L4_N2;
   wire CLK_R_M__L4_N1;
   wire CLK_R_M__L4_N0;
   wire CLK_R_M__L3_N1;
   wire CLK_R_M__L3_N0;
   wire CLK_R_M__L2_N0;
   wire CLK_R_M__L1_N0;
   wire ALU_CLK__L3_N0;
   wire ALU_CLK__L2_N0;
   wire ALU_CLK__L1_N0;
   wire CLK_UART_M__L10_N0;
   wire CLK_UART_M__L9_N0;
   wire CLK_UART_M__L8_N0;
   wire CLK_UART_M__L7_N0;
   wire CLK_UART_M__L6_N0;
   wire CLK_UART_M__L5_N1;
   wire CLK_UART_M__L5_N0;
   wire CLK_UART_M__L4_N0;
   wire CLK_UART_M__L3_N0;
   wire CLK_UART_M__L2_N0;
   wire CLK_UART_M__L1_N0;
   wire TX_CLK_M__L3_N3;
   wire TX_CLK_M__L3_N2;
   wire TX_CLK_M__L3_N1;
   wire TX_CLK_M__L3_N0;
   wire TX_CLK_M__L2_N0;
   wire TX_CLK_M__L1_N0;
   wire RX_CLK_M__L3_N0;
   wire RX_CLK_M__L2_N0;
   wire RX_CLK_M__L1_N0;
   wire FE_OFN9_SE;
   wire FE_OFN4_RST_SYNC_2_mux;
   wire FE_OFN0_RST_SYNC_1_mux;
   wire CLK_R_M;
   wire CLK_UART_M;
   wire RST_M;
   wire TX_CLK;
   wire TX_CLK_M;
   wire RX_CLK;
   wire RX_CLK_M;
   wire RST_SYNC_1;
   wire RST_SYNC_1_mux;
   wire RST_SYNC_2;
   wire RST_SYNC_2_mux;
   wire Gated_EN;
   wire ALU_CLK;
   wire WrEn_RF;
   wire RdEn_RF;
   wire RdData_valid_RF;
   wire PULSE_PG;
   wire BUSY_PG;
   wire ALU_ENABLE_in;
   wire ALU_DATA_VALID_out;
   wire FIFO_WR_INC;
   wire FIFO_FULL;
   wire FIFO_EMPTY;
   wire SYNC_data_valid_RX;
   wire SYNC_EN_OUT;
   wire n3;
   wire n8;
   wire n9;
   wire n11;
   wire n12;
   wire n13;
   wire n14;
   wire n15;
   wire n19;
   wire n20;
   wire n21;
   wire n22;
   wire n30;
   wire n31;
   wire n32;
   wire n33;
   wire n34;
   wire n35;
   wire n36;
   wire n37;
   wire n38;
   wire n39;
   wire n40;
   wire n41;
   wire n42;
   wire n43;
   wire n44;
   wire [3:0] Address_RF;
   wire [7:0] WrData_RF;
   wire [7:0] RdData_RF;
   wire [7:0] REG0_OP_A;
   wire [7:0] REG1_OP_B;
   wire [7:0] REG2_UART_config;
   wire [7:0] REG3_DIV_ratio;
   wire [7:0] div_ratio_prescale;
   wire [3:0] ALU_FUN_in;
   wire [15:0] CTRL_ALU_OUT;
   wire [7:0] FIFO_WR_DATA;
   wire [7:0] FIFO_RD_DATA;
   wire [7:0] SYNC_P_DATA_RX;
   wire [7:0] CTRL_SYNC_DATA;
endmodule

